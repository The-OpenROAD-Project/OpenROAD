module gcd (clk,
    req_rdy,
    req_val,
    reset,
    resp_rdy,
    resp_val,
    req_msg,
    resp_msg);
 input clk;
 output req_rdy;
 input req_val;
 input reset;
 input resp_rdy;
 output resp_val;
 input [31:0] req_msg;
 output [15:0] resp_msg;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire net15;
 wire net12;
 wire net14;
 wire net13;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire net11;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire net10;
 wire _143_;
 wire _144_;
 wire _145_;
 wire net9;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire net8;
 wire _158_;
 wire _159_;
 wire net7;
 wire net6;
 wire _162_;
 wire net5;
 wire _164_;
 wire net4;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire net3;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire net2;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire net1;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire \dpath.a_lt_b$in0[10] ;
 wire \dpath.a_lt_b$in0[11] ;
 wire \dpath.a_lt_b$in0[12] ;
 wire \dpath.a_lt_b$in0[13] ;
 wire \dpath.a_lt_b$in0[14] ;
 wire \dpath.a_lt_b$in0[15] ;
 wire \dpath.a_lt_b$in0[1] ;
 wire \dpath.a_lt_b$in0[2] ;
 wire \dpath.a_lt_b$in0[3] ;
 wire \dpath.a_lt_b$in0[4] ;
 wire \dpath.a_lt_b$in0[5] ;
 wire \dpath.a_lt_b$in0[6] ;
 wire \dpath.a_lt_b$in0[7] ;
 wire \dpath.a_lt_b$in0[8] ;
 wire \dpath.a_lt_b$in0[9] ;
 wire \dpath.a_lt_b$in1[0] ;
 wire \dpath.a_lt_b$in1[1] ;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net83;
 wire net82;
 wire net84;
 wire net85;
 wire clknet_2_3__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire net86;
 wire clknet_2_0__leaf_clk;
 wire clknet_0_clk;

 BUFx2_ASAP7_75t_L input15 (.A(req_msg[22]),
    .Y(net15));
 INVx1_ASAP7_75t_R _298_ (.A(_003_),
    .Y(net36));
 BUFx2_ASAP7_75t_L input14 (.A(req_msg[21]),
    .Y(net14));
 BUFx2_ASAP7_75t_L input13 (.A(req_msg[20]),
    .Y(net13));
 BUFx2_ASAP7_75t_L input12 (.A(req_msg[1]),
    .Y(net12));
 INVx1_ASAP7_75t_R _302_ (.A(_066_),
    .Y(\dpath.a_lt_b$in1[1] ));
 INVx1_ASAP7_75t_R _303_ (.A(_004_),
    .Y(\dpath.a_lt_b$in1[0] ));
 OA211x2_ASAP7_75t_SL _304_ (.A1(_052_),
    .A2(_050_),
    .B(_049_),
    .C(_046_),
    .Y(_107_));
 AO21x1_ASAP7_75t_R _305_ (.A1(_046_),
    .A2(_047_),
    .B(_044_),
    .Y(_108_));
 OA21x2_ASAP7_75t_SL _306_ (.A1(_107_),
    .A2(_108_),
    .B(_043_),
    .Y(_109_));
 OR2x2_ASAP7_75t_SL _307_ (.A(_041_),
    .B(_109_),
    .Y(_110_));
 AOI21x1_ASAP7_75t_R _308_ (.A1(_040_),
    .A2(_110_),
    .B(_038_),
    .Y(_111_));
 INVx1_ASAP7_75t_R _309_ (.A(_023_),
    .Y(_112_));
 OA21x2_ASAP7_75t_R _310_ (.A1(_065_),
    .A2(_112_),
    .B(_064_),
    .Y(_113_));
 OR3x1_ASAP7_75t_R _311_ (.A(net85),
    .B(net84),
    .C(_056_),
    .Y(_114_));
 OA21x2_ASAP7_75t_SL _312_ (.A1(net85),
    .A2(_061_),
    .B(_058_),
    .Y(_115_));
 OA21x2_ASAP7_75t_SL _313_ (.A1(_056_),
    .A2(_115_),
    .B(_055_),
    .Y(_116_));
 OA21x2_ASAP7_75t_SL _314_ (.A1(_113_),
    .A2(_114_),
    .B(_116_),
    .Y(_117_));
 OR3x1_ASAP7_75t_SL _315_ (.A(_047_),
    .B(_053_),
    .C(_050_),
    .Y(_118_));
 NOR2x1_ASAP7_75t_SL _316_ (.A(_041_),
    .B(_044_),
    .Y(_119_));
 INVx1_ASAP7_75t_R _317_ (.A(_119_),
    .Y(_120_));
 OR3x1_ASAP7_75t_L _318_ (.A(_038_),
    .B(_118_),
    .C(_120_),
    .Y(_121_));
 OAI21x1_ASAP7_75t_R _319_ (.A1(_117_),
    .A2(_121_),
    .B(_037_),
    .Y(_122_));
 OA21x2_ASAP7_75t_SL _320_ (.A1(_034_),
    .A2(_032_),
    .B(_031_),
    .Y(_123_));
 OR2x2_ASAP7_75t_SL _321_ (.A(_029_),
    .B(_123_),
    .Y(_124_));
 AO21x1_ASAP7_75t_R _322_ (.A1(_028_),
    .A2(_124_),
    .B(_026_),
    .Y(_125_));
 NAND2x1_ASAP7_75t_R _323_ (.A(_025_),
    .B(_125_),
    .Y(_126_));
 AO21x1_ASAP7_75t_SL _324_ (.A1(_034_),
    .A2(_035_),
    .B(_032_),
    .Y(_127_));
 AO21x1_ASAP7_75t_R _325_ (.A1(_031_),
    .A2(_127_),
    .B(_029_),
    .Y(_128_));
 AO21x1_ASAP7_75t_R _326_ (.A1(_028_),
    .A2(_128_),
    .B(_026_),
    .Y(_129_));
 NAND2x1_ASAP7_75t_R _327_ (.A(_025_),
    .B(_129_),
    .Y(_130_));
 OA31x2_ASAP7_75t_SL _328_ (.A1(_111_),
    .A2(_122_),
    .A3(_126_),
    .B1(_130_),
    .Y(_131_));
 BUFx2_ASAP7_75t_L input11 (.A(req_msg[19]),
    .Y(net11));
 AND4x1_ASAP7_75t_SL _330_ (.A(_042_),
    .B(_024_),
    .C(_027_),
    .D(_030_),
    .Y(_133_));
 AND5x1_ASAP7_75t_R _331_ (.A(_033_),
    .B(_036_),
    .C(_039_),
    .D(_004_),
    .E(_133_),
    .Y(_134_));
 AND4x1_ASAP7_75t_R _332_ (.A(_045_),
    .B(_048_),
    .C(_051_),
    .D(_066_),
    .Y(_135_));
 AND4x1_ASAP7_75t_R _333_ (.A(_054_),
    .B(_057_),
    .C(_060_),
    .D(_063_),
    .Y(_136_));
 AND3x1_ASAP7_75t_R _334_ (.A(_134_),
    .B(_135_),
    .C(_136_),
    .Y(_137_));
 AO21x1_ASAP7_75t_R _335_ (.A1(_131_),
    .A2(_137_),
    .B(_019_),
    .Y(_138_));
 NAND2x1_ASAP7_75t_R _336_ (.A(net33),
    .B(net86),
    .Y(_139_));
 AOI21x1_ASAP7_75t_R _337_ (.A1(_138_),
    .A2(_139_),
    .B(net34),
    .Y(_002_));
 NAND2x1_ASAP7_75t_R _338_ (.A(_003_),
    .B(_019_),
    .Y(_140_));
 NOR2x1_ASAP7_75t_R _339_ (.A(_020_),
    .B(_140_),
    .Y(net53));
 INVx1_ASAP7_75t_R _340_ (.A(net33),
    .Y(_141_));
 BUFx2_ASAP7_75t_L input10 (.A(req_msg[18]),
    .Y(net10));
 AO221x1_ASAP7_75t_SL _342_ (.A1(_141_),
    .A2(net86),
    .B1(net53),
    .B2(net35),
    .C(net34),
    .Y(_000_));
 INVx1_ASAP7_75t_R _343_ (.A(_019_),
    .Y(_143_));
 AND3x1_ASAP7_75t_R _344_ (.A(_143_),
    .B(_131_),
    .C(_137_),
    .Y(_144_));
 AND2x2_ASAP7_75t_SL _345_ (.A(_003_),
    .B(_019_),
    .Y(_145_));
 BUFx2_ASAP7_75t_L input9 (.A(req_msg[17]),
    .Y(net9));
 AOI21x1_ASAP7_75t_R _347_ (.A1(net35),
    .A2(_145_),
    .B(_020_),
    .Y(_147_));
 INVx1_ASAP7_75t_R _348_ (.A(net34),
    .Y(_148_));
 OA21x2_ASAP7_75t_SL _349_ (.A1(_144_),
    .A2(_147_),
    .B(_148_),
    .Y(_001_));
 INVx1_ASAP7_75t_R _350_ (.A(_005_),
    .Y(\dpath.a_lt_b$in0[9] ));
 INVx1_ASAP7_75t_R _351_ (.A(_006_),
    .Y(\dpath.a_lt_b$in0[8] ));
 INVx1_ASAP7_75t_R _352_ (.A(_007_),
    .Y(\dpath.a_lt_b$in0[7] ));
 INVx1_ASAP7_75t_R _353_ (.A(_008_),
    .Y(\dpath.a_lt_b$in0[6] ));
 INVx1_ASAP7_75t_R _354_ (.A(_009_),
    .Y(\dpath.a_lt_b$in0[5] ));
 INVx1_ASAP7_75t_R _355_ (.A(_010_),
    .Y(\dpath.a_lt_b$in0[4] ));
 INVx1_ASAP7_75t_R _356_ (.A(_011_),
    .Y(\dpath.a_lt_b$in0[3] ));
 INVx1_ASAP7_75t_R _357_ (.A(_012_),
    .Y(\dpath.a_lt_b$in0[2] ));
 INVx1_ASAP7_75t_R _358_ (.A(_022_),
    .Y(\dpath.a_lt_b$in0[1] ));
 INVx1_ASAP7_75t_R _359_ (.A(_013_),
    .Y(\dpath.a_lt_b$in0[15] ));
 INVx1_ASAP7_75t_R _360_ (.A(_014_),
    .Y(\dpath.a_lt_b$in0[14] ));
 INVx1_ASAP7_75t_R _361_ (.A(_015_),
    .Y(\dpath.a_lt_b$in0[13] ));
 INVx1_ASAP7_75t_R _362_ (.A(_016_),
    .Y(\dpath.a_lt_b$in0[12] ));
 INVx1_ASAP7_75t_R _363_ (.A(_017_),
    .Y(\dpath.a_lt_b$in0[11] ));
 INVx1_ASAP7_75t_R _364_ (.A(_018_),
    .Y(\dpath.a_lt_b$in0[10] ));
 AND2x2_ASAP7_75t_R _365_ (.A(_003_),
    .B(_143_),
    .Y(_149_));
 AND2x2_ASAP7_75t_R _366_ (.A(_131_),
    .B(_149_),
    .Y(_150_));
 NAND2x1_ASAP7_75t_R _367_ (.A(net37),
    .B(_150_),
    .Y(_151_));
 AO21x1_ASAP7_75t_SL _368_ (.A1(_040_),
    .A2(_110_),
    .B(_038_),
    .Y(_152_));
 OA21x2_ASAP7_75t_SL _369_ (.A1(_117_),
    .A2(_121_),
    .B(_037_),
    .Y(_153_));
 AND3x1_ASAP7_75t_SL _370_ (.A(_152_),
    .B(_153_),
    .C(_125_),
    .Y(_154_));
 AND3x1_ASAP7_75t_R _371_ (.A(_025_),
    .B(_003_),
    .C(_143_),
    .Y(_155_));
 OAI21x1_ASAP7_75t_SL _372_ (.A1(_154_),
    .A2(_129_),
    .B(_155_),
    .Y(_156_));
 BUFx2_ASAP7_75t_L input8 (.A(req_msg[16]),
    .Y(net8));
 NAND2x1_ASAP7_75t_R _374_ (.A(net86),
    .B(net8),
    .Y(_158_));
 OA211x2_ASAP7_75t_SL _375_ (.A1(_004_),
    .A2(net83),
    .B(_158_),
    .C(_140_),
    .Y(_159_));
 AOI22x1_ASAP7_75t_SL _376_ (.A1(_070_),
    .A2(_145_),
    .B1(_151_),
    .B2(_159_),
    .Y(_071_));
 BUFx2_ASAP7_75t_L input7 (.A(req_msg[15]),
    .Y(net7));
 BUFx2_ASAP7_75t_L input6 (.A(req_msg[14]),
    .Y(net6));
 NOR2x1_ASAP7_75t_R _379_ (.A(_039_),
    .B(net83),
    .Y(_162_));
 BUFx2_ASAP7_75t_L input5 (.A(req_msg[13]),
    .Y(net5));
 AO21x1_ASAP7_75t_R _381_ (.A1(net86),
    .A2(net19),
    .B(_145_),
    .Y(_164_));
 BUFx2_ASAP7_75t_L input4 (.A(req_msg[12]),
    .Y(net4));
 OR2x2_ASAP7_75t_R _383_ (.A(_044_),
    .B(_118_),
    .Y(_166_));
 OA21x2_ASAP7_75t_SL _384_ (.A1(_117_),
    .A2(_166_),
    .B(_109_),
    .Y(_167_));
 XOR2x2_ASAP7_75t_R _385_ (.A(_041_),
    .B(_167_),
    .Y(net38));
 AND3x1_ASAP7_75t_R _386_ (.A(_131_),
    .B(_149_),
    .C(net38),
    .Y(_168_));
 OA33x2_ASAP7_75t_SL _387_ (.A1(net86),
    .A2(\dpath.a_lt_b$in0[10] ),
    .A3(_143_),
    .B1(_162_),
    .B2(_164_),
    .B3(_168_),
    .Y(_072_));
 NAND2x1_ASAP7_75t_R _388_ (.A(net86),
    .B(net20),
    .Y(_169_));
 OA211x2_ASAP7_75t_SL _389_ (.A1(_036_),
    .A2(net82),
    .B(_169_),
    .C(_140_),
    .Y(_170_));
 OA21x2_ASAP7_75t_R _390_ (.A1(_041_),
    .A2(_043_),
    .B(_040_),
    .Y(_171_));
 INVx3_ASAP7_75t_SL _391_ (.A(_069_),
    .Y(_021_));
 OA21x2_ASAP7_75t_R _392_ (.A1(_021_),
    .A2(_068_),
    .B(_067_),
    .Y(_172_));
 OR3x1_ASAP7_75t_R _393_ (.A(net85),
    .B(net84),
    .C(_065_),
    .Y(_173_));
 OR3x1_ASAP7_75t_L _394_ (.A(net85),
    .B(_064_),
    .C(net84),
    .Y(_174_));
 OA211x2_ASAP7_75t_SL _395_ (.A1(_172_),
    .A2(_173_),
    .B(_115_),
    .C(_174_),
    .Y(_175_));
 OR2x2_ASAP7_75t_R _396_ (.A(_056_),
    .B(_118_),
    .Y(_176_));
 OR2x2_ASAP7_75t_R _397_ (.A(_053_),
    .B(_055_),
    .Y(_177_));
 OR2x2_ASAP7_75t_R _398_ (.A(_047_),
    .B(_050_),
    .Y(_178_));
 AO21x1_ASAP7_75t_R _399_ (.A1(_052_),
    .A2(_177_),
    .B(_178_),
    .Y(_179_));
 OA21x2_ASAP7_75t_SL _400_ (.A1(_175_),
    .A2(_176_),
    .B(_179_),
    .Y(_180_));
 OA21x2_ASAP7_75t_R _401_ (.A1(_047_),
    .A2(_049_),
    .B(_046_),
    .Y(_181_));
 AO21x2_ASAP7_75t_SL _402_ (.A1(_180_),
    .A2(_181_),
    .B(_120_),
    .Y(_182_));
 INVx1_ASAP7_75t_R _403_ (.A(_038_),
    .Y(_183_));
 AO21x1_ASAP7_75t_R _404_ (.A1(_171_),
    .A2(_182_),
    .B(_183_),
    .Y(_184_));
 NAND3x1_ASAP7_75t_R _405_ (.A(_183_),
    .B(_171_),
    .C(_182_),
    .Y(_185_));
 NAND2x1_ASAP7_75t_R _406_ (.A(_131_),
    .B(_149_),
    .Y(_186_));
 AO21x1_ASAP7_75t_R _407_ (.A1(_184_),
    .A2(_185_),
    .B(_186_),
    .Y(_187_));
 AOI22x1_ASAP7_75t_SL _408_ (.A1(_017_),
    .A2(_145_),
    .B1(_170_),
    .B2(_187_),
    .Y(_073_));
 OR2x2_ASAP7_75t_R _409_ (.A(_003_),
    .B(net21),
    .Y(_188_));
 NAND2x1_ASAP7_75t_R _410_ (.A(_016_),
    .B(_145_),
    .Y(_189_));
 OAI21x1_ASAP7_75t_R _411_ (.A1(_033_),
    .A2(_131_),
    .B(_149_),
    .Y(_190_));
 NAND2x1_ASAP7_75t_R _412_ (.A(_152_),
    .B(_153_),
    .Y(_191_));
 XNOR2x2_ASAP7_75t_R _413_ (.A(_035_),
    .B(_191_),
    .Y(net40));
 AO32x1_ASAP7_75t_SL _414_ (.A1(_188_),
    .A2(_189_),
    .A3(_190_),
    .B1(net40),
    .B2(_150_),
    .Y(_074_));
 OA21x2_ASAP7_75t_R _415_ (.A1(_035_),
    .A2(_037_),
    .B(_034_),
    .Y(_192_));
 AO21x1_ASAP7_75t_R _416_ (.A1(_038_),
    .A2(_037_),
    .B(_035_),
    .Y(_193_));
 AO32x1_ASAP7_75t_SL _417_ (.A1(_171_),
    .A2(_182_),
    .A3(_192_),
    .B1(_193_),
    .B2(_034_),
    .Y(_194_));
 XOR2x2_ASAP7_75t_SL _418_ (.A(_032_),
    .B(_194_),
    .Y(net41));
 BUFx2_ASAP7_75t_L input3 (.A(req_msg[11]),
    .Y(net3));
 AOI21x1_ASAP7_75t_R _420_ (.A1(net86),
    .A2(net22),
    .B(_145_),
    .Y(_196_));
 OAI21x1_ASAP7_75t_R _421_ (.A1(_030_),
    .A2(net82),
    .B(_196_),
    .Y(_197_));
 NAND2x1_ASAP7_75t_R _422_ (.A(_015_),
    .B(_145_),
    .Y(_198_));
 AO32x1_ASAP7_75t_SL _423_ (.A1(_131_),
    .A2(_149_),
    .A3(net41),
    .B1(_197_),
    .B2(_198_),
    .Y(_075_));
 OR2x2_ASAP7_75t_R _424_ (.A(_003_),
    .B(net24),
    .Y(_199_));
 NAND2x1_ASAP7_75t_R _425_ (.A(_014_),
    .B(_145_),
    .Y(_200_));
 OAI21x1_ASAP7_75t_R _426_ (.A1(_027_),
    .A2(_131_),
    .B(_149_),
    .Y(_201_));
 AO32x1_ASAP7_75t_R _427_ (.A1(_152_),
    .A2(_153_),
    .A3(_123_),
    .B1(_127_),
    .B2(_031_),
    .Y(_202_));
 XOR2x2_ASAP7_75t_SL _428_ (.A(_029_),
    .B(_202_),
    .Y(net42));
 AO32x1_ASAP7_75t_SL _429_ (.A1(_199_),
    .A2(_200_),
    .A3(_201_),
    .B1(net42),
    .B2(_150_),
    .Y(_076_));
 OA21x2_ASAP7_75t_R _430_ (.A1(_032_),
    .A2(_192_),
    .B(_031_),
    .Y(_203_));
 OA21x2_ASAP7_75t_R _431_ (.A1(_029_),
    .A2(_203_),
    .B(_171_),
    .Y(_204_));
 AND3x1_ASAP7_75t_SL _432_ (.A(_180_),
    .B(_181_),
    .C(_204_),
    .Y(_205_));
 AO21x1_ASAP7_75t_R _433_ (.A1(_034_),
    .A2(_193_),
    .B(_032_),
    .Y(_206_));
 AND2x2_ASAP7_75t_R _434_ (.A(_120_),
    .B(_171_),
    .Y(_207_));
 AO221x1_ASAP7_75t_R _435_ (.A1(_031_),
    .A2(_206_),
    .B1(_207_),
    .B2(_203_),
    .C(_029_),
    .Y(_208_));
 OA21x2_ASAP7_75t_R _436_ (.A1(_205_),
    .A2(_208_),
    .B(_028_),
    .Y(_209_));
 XOR2x2_ASAP7_75t_SL _437_ (.A(_026_),
    .B(_209_),
    .Y(net43));
 NAND2x1_ASAP7_75t_R _438_ (.A(_013_),
    .B(_145_),
    .Y(_210_));
 OAI21x1_ASAP7_75t_R _439_ (.A1(_024_),
    .A2(_131_),
    .B(_149_),
    .Y(_211_));
 OA211x2_ASAP7_75t_R _440_ (.A1(_003_),
    .A2(net25),
    .B(_210_),
    .C(_211_),
    .Y(_212_));
 AO21x1_ASAP7_75t_SL _441_ (.A1(_150_),
    .A2(net43),
    .B(_212_),
    .Y(_077_));
 AND3x1_ASAP7_75t_R _442_ (.A(net44),
    .B(_131_),
    .C(_149_),
    .Y(_213_));
 AO21x1_ASAP7_75t_R _443_ (.A1(net86),
    .A2(net9),
    .B(_145_),
    .Y(_214_));
 BUFx2_ASAP7_75t_L input2 (.A(req_msg[10]),
    .Y(net2));
 NOR2x1_ASAP7_75t_SL _445_ (.A(_066_),
    .B(net83),
    .Y(_216_));
 OA33x2_ASAP7_75t_SL _446_ (.A1(net86),
    .A2(\dpath.a_lt_b$in0[1] ),
    .A3(_143_),
    .B1(_213_),
    .B2(_214_),
    .B3(_216_),
    .Y(_078_));
 XNOR2x2_ASAP7_75t_R _447_ (.A(_065_),
    .B(_023_),
    .Y(net45));
 AND3x1_ASAP7_75t_SL _448_ (.A(_131_),
    .B(_149_),
    .C(net45),
    .Y(_217_));
 AO21x1_ASAP7_75t_R _449_ (.A1(net86),
    .A2(net10),
    .B(_145_),
    .Y(_218_));
 NOR2x1_ASAP7_75t_SL _450_ (.A(_063_),
    .B(net83),
    .Y(_219_));
 OA33x2_ASAP7_75t_SL _451_ (.A1(net86),
    .A2(\dpath.a_lt_b$in0[2] ),
    .A3(_143_),
    .B1(_217_),
    .B2(_218_),
    .B3(_219_),
    .Y(_079_));
 OA21x2_ASAP7_75t_R _452_ (.A1(_065_),
    .A2(_172_),
    .B(_064_),
    .Y(_220_));
 XOR2x2_ASAP7_75t_R _453_ (.A(net84),
    .B(_220_),
    .Y(net46));
 AND3x1_ASAP7_75t_SL _454_ (.A(_131_),
    .B(_149_),
    .C(net46),
    .Y(_221_));
 AO21x1_ASAP7_75t_R _455_ (.A1(net86),
    .A2(net11),
    .B(_145_),
    .Y(_222_));
 NOR2x1_ASAP7_75t_SL _456_ (.A(_060_),
    .B(net83),
    .Y(_223_));
 OA33x2_ASAP7_75t_SL _457_ (.A1(net86),
    .A2(\dpath.a_lt_b$in0[3] ),
    .A3(_143_),
    .B1(_221_),
    .B2(_222_),
    .B3(_223_),
    .Y(_080_));
 OA21x2_ASAP7_75t_R _458_ (.A1(net84),
    .A2(_113_),
    .B(_061_),
    .Y(_224_));
 XOR2x2_ASAP7_75t_R _459_ (.A(net85),
    .B(_224_),
    .Y(net47));
 AND3x1_ASAP7_75t_R _460_ (.A(_131_),
    .B(_149_),
    .C(net47),
    .Y(_225_));
 AO21x1_ASAP7_75t_R _461_ (.A1(net86),
    .A2(net13),
    .B(_145_),
    .Y(_226_));
 NOR2x1_ASAP7_75t_SL _462_ (.A(_057_),
    .B(net83),
    .Y(_227_));
 OA33x2_ASAP7_75t_SL _463_ (.A1(net86),
    .A2(\dpath.a_lt_b$in0[4] ),
    .A3(_143_),
    .B1(_225_),
    .B2(_226_),
    .B3(_227_),
    .Y(_081_));
 XOR2x2_ASAP7_75t_R _464_ (.A(_056_),
    .B(_175_),
    .Y(net48));
 AND3x1_ASAP7_75t_R _465_ (.A(_131_),
    .B(_149_),
    .C(net48),
    .Y(_228_));
 AO21x1_ASAP7_75t_R _466_ (.A1(net86),
    .A2(net14),
    .B(_145_),
    .Y(_229_));
 NOR2x1_ASAP7_75t_SL _467_ (.A(_054_),
    .B(net83),
    .Y(_230_));
 OA33x2_ASAP7_75t_SL _468_ (.A1(net86),
    .A2(\dpath.a_lt_b$in0[5] ),
    .A3(_143_),
    .B1(_228_),
    .B2(_229_),
    .B3(_230_),
    .Y(_082_));
 XOR2x2_ASAP7_75t_R _469_ (.A(_053_),
    .B(_117_),
    .Y(net49));
 AND3x1_ASAP7_75t_R _470_ (.A(_131_),
    .B(_149_),
    .C(net49),
    .Y(_231_));
 AO21x1_ASAP7_75t_R _471_ (.A1(net86),
    .A2(net15),
    .B(_145_),
    .Y(_232_));
 NOR2x1_ASAP7_75t_SL _472_ (.A(_051_),
    .B(net83),
    .Y(_233_));
 OA33x2_ASAP7_75t_SL _473_ (.A1(net86),
    .A2(\dpath.a_lt_b$in0[6] ),
    .A3(_143_),
    .B1(_231_),
    .B2(_232_),
    .B3(_233_),
    .Y(_083_));
 OR3x1_ASAP7_75t_SL _474_ (.A(_053_),
    .B(_056_),
    .C(_175_),
    .Y(_234_));
 AND3x1_ASAP7_75t_SL _475_ (.A(_052_),
    .B(_177_),
    .C(_234_),
    .Y(_235_));
 XOR2x2_ASAP7_75t_R _476_ (.A(_050_),
    .B(_235_),
    .Y(net50));
 AND2x2_ASAP7_75t_SL _477_ (.A(_150_),
    .B(net50),
    .Y(_236_));
 AO21x1_ASAP7_75t_R _478_ (.A1(net86),
    .A2(net16),
    .B(_145_),
    .Y(_237_));
 NOR2x1_ASAP7_75t_R _479_ (.A(_048_),
    .B(net83),
    .Y(_238_));
 OA33x2_ASAP7_75t_SL _480_ (.A1(net86),
    .A2(\dpath.a_lt_b$in0[7] ),
    .A3(_143_),
    .B1(_236_),
    .B2(_237_),
    .B3(_238_),
    .Y(_084_));
 NOR2x1_ASAP7_75t_SL _481_ (.A(_045_),
    .B(net83),
    .Y(_239_));
 AO21x1_ASAP7_75t_R _482_ (.A1(net86),
    .A2(net17),
    .B(_145_),
    .Y(_240_));
 OA21x2_ASAP7_75t_SL _483_ (.A1(_053_),
    .A2(_117_),
    .B(_052_),
    .Y(_241_));
 OA21x2_ASAP7_75t_SL _484_ (.A1(_050_),
    .A2(_241_),
    .B(_049_),
    .Y(_242_));
 XOR2x2_ASAP7_75t_L _485_ (.A(_047_),
    .B(_242_),
    .Y(net51));
 AND3x1_ASAP7_75t_SL _486_ (.A(_131_),
    .B(_149_),
    .C(net51),
    .Y(_243_));
 OA33x2_ASAP7_75t_SL _487_ (.A1(net86),
    .A2(\dpath.a_lt_b$in0[8] ),
    .A3(_143_),
    .B1(_239_),
    .B2(_240_),
    .B3(_243_),
    .Y(_085_));
 NOR2x1_ASAP7_75t_R _488_ (.A(_042_),
    .B(net83),
    .Y(_244_));
 AO21x1_ASAP7_75t_R _489_ (.A1(net86),
    .A2(net18),
    .B(_145_),
    .Y(_245_));
 NAND2x1_ASAP7_75t_R _490_ (.A(_180_),
    .B(_181_),
    .Y(_246_));
 XNOR2x2_ASAP7_75t_R _491_ (.A(_044_),
    .B(_246_),
    .Y(net52));
 AND2x2_ASAP7_75t_SL _492_ (.A(_150_),
    .B(net52),
    .Y(_247_));
 OA33x2_ASAP7_75t_SL _493_ (.A1(net86),
    .A2(\dpath.a_lt_b$in0[9] ),
    .A3(_143_),
    .B1(_244_),
    .B2(_245_),
    .B3(_247_),
    .Y(_086_));
 BUFx2_ASAP7_75t_L input1 (.A(req_msg[0]),
    .Y(net1));
 AND2x2_ASAP7_75t_R _495_ (.A(_003_),
    .B(\dpath.a_lt_b$in1[0] ),
    .Y(_249_));
 AO21x1_ASAP7_75t_R _496_ (.A1(net86),
    .A2(net1),
    .B(_249_),
    .Y(_250_));
 NOR2x1_ASAP7_75t_R _497_ (.A(_070_),
    .B(net83),
    .Y(_251_));
 AO21x1_ASAP7_75t_SL _498_ (.A1(net83),
    .A2(_250_),
    .B(_251_),
    .Y(_087_));
 NOR2x1_ASAP7_75t_R _499_ (.A(\dpath.a_lt_b$in0[10] ),
    .B(net83),
    .Y(_252_));
 NAND2x1_ASAP7_75t_R _500_ (.A(net86),
    .B(net2),
    .Y(_253_));
 OA211x2_ASAP7_75t_SL _501_ (.A1(net86),
    .A2(_039_),
    .B(net83),
    .C(_253_),
    .Y(_254_));
 NOR2x2_ASAP7_75t_SL _502_ (.A(_252_),
    .B(_254_),
    .Y(_088_));
 NOR2x1_ASAP7_75t_R _503_ (.A(\dpath.a_lt_b$in0[11] ),
    .B(net82),
    .Y(_255_));
 NAND2x1_ASAP7_75t_R _504_ (.A(net86),
    .B(net3),
    .Y(_256_));
 OA211x2_ASAP7_75t_SL _505_ (.A1(net86),
    .A2(_036_),
    .B(net82),
    .C(_256_),
    .Y(_257_));
 NOR2x2_ASAP7_75t_SL _506_ (.A(_255_),
    .B(_257_),
    .Y(_089_));
 NOR2x1_ASAP7_75t_R _507_ (.A(\dpath.a_lt_b$in0[12] ),
    .B(net82),
    .Y(_258_));
 NAND2x1_ASAP7_75t_R _508_ (.A(net86),
    .B(net4),
    .Y(_259_));
 OA211x2_ASAP7_75t_SL _509_ (.A1(net86),
    .A2(_033_),
    .B(net82),
    .C(_259_),
    .Y(_260_));
 NOR2x2_ASAP7_75t_SL _510_ (.A(_258_),
    .B(_260_),
    .Y(_090_));
 NOR2x1_ASAP7_75t_R _511_ (.A(\dpath.a_lt_b$in0[13] ),
    .B(net82),
    .Y(_261_));
 NAND2x1_ASAP7_75t_R _512_ (.A(net86),
    .B(net5),
    .Y(_262_));
 OA211x2_ASAP7_75t_SL _513_ (.A1(net86),
    .A2(_030_),
    .B(net82),
    .C(_262_),
    .Y(_263_));
 NOR2x2_ASAP7_75t_SL _514_ (.A(_261_),
    .B(_263_),
    .Y(_091_));
 NOR2x1_ASAP7_75t_R _515_ (.A(\dpath.a_lt_b$in0[14] ),
    .B(net82),
    .Y(_264_));
 NAND2x1_ASAP7_75t_R _516_ (.A(net86),
    .B(net6),
    .Y(_265_));
 OA211x2_ASAP7_75t_SL _517_ (.A1(net86),
    .A2(_027_),
    .B(net82),
    .C(_265_),
    .Y(_266_));
 NOR2x2_ASAP7_75t_SL _518_ (.A(_264_),
    .B(_266_),
    .Y(_092_));
 NOR2x1_ASAP7_75t_R _519_ (.A(\dpath.a_lt_b$in0[15] ),
    .B(net82),
    .Y(_267_));
 NAND2x1_ASAP7_75t_R _520_ (.A(net86),
    .B(net7),
    .Y(_268_));
 OA211x2_ASAP7_75t_SL _521_ (.A1(net86),
    .A2(_024_),
    .B(net82),
    .C(_268_),
    .Y(_269_));
 NOR2x2_ASAP7_75t_SL _522_ (.A(_267_),
    .B(_269_),
    .Y(_093_));
 AND2x2_ASAP7_75t_R _523_ (.A(_003_),
    .B(\dpath.a_lt_b$in1[1] ),
    .Y(_270_));
 AO21x1_ASAP7_75t_R _524_ (.A1(net86),
    .A2(net12),
    .B(_270_),
    .Y(_271_));
 NOR2x1_ASAP7_75t_R _525_ (.A(_022_),
    .B(net83),
    .Y(_272_));
 AO21x1_ASAP7_75t_SL _526_ (.A1(net83),
    .A2(_271_),
    .B(_272_),
    .Y(_094_));
 NOR2x1_ASAP7_75t_R _527_ (.A(\dpath.a_lt_b$in0[2] ),
    .B(net83),
    .Y(_273_));
 NAND2x1_ASAP7_75t_R _528_ (.A(net86),
    .B(net23),
    .Y(_274_));
 OA211x2_ASAP7_75t_SL _529_ (.A1(net86),
    .A2(_063_),
    .B(net83),
    .C(_274_),
    .Y(_275_));
 NOR2x2_ASAP7_75t_SL _530_ (.A(_273_),
    .B(_275_),
    .Y(_095_));
 NOR2x1_ASAP7_75t_R _531_ (.A(\dpath.a_lt_b$in0[3] ),
    .B(net83),
    .Y(_276_));
 NAND2x1_ASAP7_75t_R _532_ (.A(net86),
    .B(net26),
    .Y(_277_));
 OA211x2_ASAP7_75t_SL _533_ (.A1(net86),
    .A2(_060_),
    .B(net83),
    .C(_277_),
    .Y(_278_));
 NOR2x2_ASAP7_75t_SL _534_ (.A(_276_),
    .B(_278_),
    .Y(_096_));
 NOR2x1_ASAP7_75t_R _535_ (.A(\dpath.a_lt_b$in0[4] ),
    .B(net83),
    .Y(_279_));
 NAND2x1_ASAP7_75t_R _536_ (.A(net86),
    .B(net27),
    .Y(_280_));
 OA211x2_ASAP7_75t_SL _537_ (.A1(net86),
    .A2(_057_),
    .B(net83),
    .C(_280_),
    .Y(_281_));
 NOR2x2_ASAP7_75t_SL _538_ (.A(_279_),
    .B(_281_),
    .Y(_097_));
 NOR2x1_ASAP7_75t_R _539_ (.A(\dpath.a_lt_b$in0[5] ),
    .B(net83),
    .Y(_282_));
 NAND2x1_ASAP7_75t_R _540_ (.A(net86),
    .B(net28),
    .Y(_283_));
 OA211x2_ASAP7_75t_R _541_ (.A1(net86),
    .A2(_054_),
    .B(net83),
    .C(_283_),
    .Y(_284_));
 NOR2x1_ASAP7_75t_SL _542_ (.A(_282_),
    .B(_284_),
    .Y(_098_));
 NOR2x1_ASAP7_75t_R _543_ (.A(\dpath.a_lt_b$in0[6] ),
    .B(net83),
    .Y(_285_));
 NAND2x1_ASAP7_75t_R _544_ (.A(net86),
    .B(net29),
    .Y(_286_));
 OA211x2_ASAP7_75t_R _545_ (.A1(net86),
    .A2(_051_),
    .B(net83),
    .C(_286_),
    .Y(_287_));
 NOR2x1_ASAP7_75t_SL _546_ (.A(_285_),
    .B(_287_),
    .Y(_099_));
 NOR2x1_ASAP7_75t_R _547_ (.A(\dpath.a_lt_b$in0[7] ),
    .B(net83),
    .Y(_288_));
 NAND2x1_ASAP7_75t_R _548_ (.A(net86),
    .B(net30),
    .Y(_289_));
 OA211x2_ASAP7_75t_R _549_ (.A1(net86),
    .A2(_048_),
    .B(net83),
    .C(_289_),
    .Y(_290_));
 NOR2x1_ASAP7_75t_SL _550_ (.A(_288_),
    .B(_290_),
    .Y(_100_));
 NOR2x1_ASAP7_75t_R _551_ (.A(\dpath.a_lt_b$in0[8] ),
    .B(net83),
    .Y(_291_));
 NAND2x1_ASAP7_75t_R _552_ (.A(net86),
    .B(net31),
    .Y(_292_));
 OA211x2_ASAP7_75t_R _553_ (.A1(net86),
    .A2(_045_),
    .B(net83),
    .C(_292_),
    .Y(_293_));
 NOR2x1_ASAP7_75t_SL _554_ (.A(_291_),
    .B(_293_),
    .Y(_101_));
 NOR2x1_ASAP7_75t_R _555_ (.A(\dpath.a_lt_b$in0[9] ),
    .B(net83),
    .Y(_294_));
 NAND2x1_ASAP7_75t_R _556_ (.A(net86),
    .B(net32),
    .Y(_295_));
 OA211x2_ASAP7_75t_R _557_ (.A1(net86),
    .A2(_042_),
    .B(net83),
    .C(_295_),
    .Y(_296_));
 NOR2x1_ASAP7_75t_SL _558_ (.A(_294_),
    .B(_296_),
    .Y(_102_));
 NAND2x1_ASAP7_75t_R _559_ (.A(_184_),
    .B(_185_),
    .Y(net39));
 FAx1_ASAP7_75t_R _560_ (.SN(net44),
    .A(_021_),
    .B(\dpath.a_lt_b$in1[1] ),
    .CI(_022_),
    .CON(_023_));
 HAxp5_ASAP7_75t_R _561_ (.A(_024_),
    .B(\dpath.a_lt_b$in0[15] ),
    .CON(_025_),
    .SN(_026_));
 HAxp5_ASAP7_75t_R _562_ (.A(_027_),
    .B(\dpath.a_lt_b$in0[14] ),
    .CON(_028_),
    .SN(_029_));
 HAxp5_ASAP7_75t_R _563_ (.A(_030_),
    .B(\dpath.a_lt_b$in0[13] ),
    .CON(_031_),
    .SN(_032_));
 HAxp5_ASAP7_75t_R _564_ (.A(_033_),
    .B(\dpath.a_lt_b$in0[12] ),
    .CON(_034_),
    .SN(_035_));
 HAxp5_ASAP7_75t_R _565_ (.A(_036_),
    .B(\dpath.a_lt_b$in0[11] ),
    .CON(_037_),
    .SN(_038_));
 HAxp5_ASAP7_75t_R _566_ (.A(_039_),
    .B(\dpath.a_lt_b$in0[10] ),
    .CON(_040_),
    .SN(_041_));
 HAxp5_ASAP7_75t_R _567_ (.A(_042_),
    .B(\dpath.a_lt_b$in0[9] ),
    .CON(_043_),
    .SN(_044_));
 HAxp5_ASAP7_75t_R _568_ (.A(_045_),
    .B(\dpath.a_lt_b$in0[8] ),
    .CON(_046_),
    .SN(_047_));
 HAxp5_ASAP7_75t_R _569_ (.A(_048_),
    .B(\dpath.a_lt_b$in0[7] ),
    .CON(_049_),
    .SN(_050_));
 HAxp5_ASAP7_75t_R _570_ (.A(_051_),
    .B(\dpath.a_lt_b$in0[6] ),
    .CON(_052_),
    .SN(_053_));
 HAxp5_ASAP7_75t_R _571_ (.A(_054_),
    .B(\dpath.a_lt_b$in0[5] ),
    .CON(_055_),
    .SN(_056_));
 HAxp5_ASAP7_75t_R _572_ (.A(_057_),
    .B(\dpath.a_lt_b$in0[4] ),
    .CON(_058_),
    .SN(_059_));
 HAxp5_ASAP7_75t_R _573_ (.A(_060_),
    .B(\dpath.a_lt_b$in0[3] ),
    .CON(_061_),
    .SN(_062_));
 HAxp5_ASAP7_75t_R _574_ (.A(_063_),
    .B(\dpath.a_lt_b$in0[2] ),
    .CON(_064_),
    .SN(_065_));
 HAxp5_ASAP7_75t_R _575_ (.A(_066_),
    .B(\dpath.a_lt_b$in0[1] ),
    .CON(_067_),
    .SN(_068_));
 HAxp5_ASAP7_75t_R _576_ (.A(\dpath.a_lt_b$in1[0] ),
    .B(_070_),
    .CON(_069_),
    .SN(net37));
 DFFHQNx1_ASAP7_75t_SL \ctrl.state.out[0]$_DFF_P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_000_),
    .QN(_003_));
 DFFHQNx1_ASAP7_75t_SL \ctrl.state.out[1]$_DFF_P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_001_),
    .QN(_020_));
 DFFHQNx1_ASAP7_75t_SL \ctrl.state.out[2]$_DFF_P_  (.CLK(clknet_2_3__leaf_clk),
    .D(_002_),
    .QN(_019_));
 DFFHQNx1_ASAP7_75t_SL \dpath.a_reg.out[0]$_DFFE_PP_  (.CLK(clknet_2_3__leaf_clk),
    .D(_071_),
    .QN(_070_));
 DFFHQNx1_ASAP7_75t_SL \dpath.a_reg.out[10]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .D(_072_),
    .QN(_018_));
 DFFHQNx1_ASAP7_75t_SL \dpath.a_reg.out[11]$_DFFE_PP_  (.CLK(clknet_2_3__leaf_clk),
    .D(_073_),
    .QN(_017_));
 DFFHQNx1_ASAP7_75t_SL \dpath.a_reg.out[12]$_DFFE_PP_  (.CLK(clknet_2_3__leaf_clk),
    .D(_074_),
    .QN(_016_));
 DFFHQNx1_ASAP7_75t_SL \dpath.a_reg.out[13]$_DFFE_PP_  (.CLK(clknet_2_3__leaf_clk),
    .D(_075_),
    .QN(_015_));
 DFFHQNx1_ASAP7_75t_SL \dpath.a_reg.out[14]$_DFFE_PP_  (.CLK(clknet_2_2__leaf_clk),
    .D(_076_),
    .QN(_014_));
 DFFHQNx1_ASAP7_75t_SL \dpath.a_reg.out[15]$_DFFE_PP_  (.CLK(clknet_2_2__leaf_clk),
    .D(_077_),
    .QN(_013_));
 DFFHQNx1_ASAP7_75t_SL \dpath.a_reg.out[1]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .D(_078_),
    .QN(_022_));
 DFFHQNx1_ASAP7_75t_SL \dpath.a_reg.out[2]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .D(_079_),
    .QN(_012_));
 DFFHQNx1_ASAP7_75t_SL \dpath.a_reg.out[3]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .D(_080_),
    .QN(_011_));
 DFFHQNx1_ASAP7_75t_SL \dpath.a_reg.out[4]$_DFFE_PP_  (.CLK(clknet_2_0__leaf_clk),
    .D(_081_),
    .QN(_010_));
 DFFHQNx1_ASAP7_75t_SL \dpath.a_reg.out[5]$_DFFE_PP_  (.CLK(clknet_2_0__leaf_clk),
    .D(_082_),
    .QN(_009_));
 DFFHQNx1_ASAP7_75t_SL \dpath.a_reg.out[6]$_DFFE_PP_  (.CLK(clknet_2_0__leaf_clk),
    .D(_083_),
    .QN(_008_));
 DFFHQNx1_ASAP7_75t_SL \dpath.a_reg.out[7]$_DFFE_PP_  (.CLK(clknet_2_0__leaf_clk),
    .D(_084_),
    .QN(_007_));
 DFFHQNx1_ASAP7_75t_SL \dpath.a_reg.out[8]$_DFFE_PP_  (.CLK(clknet_2_0__leaf_clk),
    .D(_085_),
    .QN(_006_));
 DFFHQNx1_ASAP7_75t_SL \dpath.a_reg.out[9]$_DFFE_PP_  (.CLK(clknet_2_2__leaf_clk),
    .D(_086_),
    .QN(_005_));
 DFFHQNx1_ASAP7_75t_SL \dpath.b_reg.out[0]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .D(_087_),
    .QN(_004_));
 DFFHQNx1_ASAP7_75t_SL \dpath.b_reg.out[10]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .D(_088_),
    .QN(_039_));
 DFFHQNx1_ASAP7_75t_SL \dpath.b_reg.out[11]$_DFFE_PP_  (.CLK(clknet_2_3__leaf_clk),
    .D(_089_),
    .QN(_036_));
 DFFHQNx1_ASAP7_75t_SL \dpath.b_reg.out[12]$_DFFE_PP_  (.CLK(clknet_2_3__leaf_clk),
    .D(_090_),
    .QN(_033_));
 DFFHQNx1_ASAP7_75t_SL \dpath.b_reg.out[13]$_DFFE_PP_  (.CLK(clknet_2_2__leaf_clk),
    .D(_091_),
    .QN(_030_));
 DFFHQNx1_ASAP7_75t_SL \dpath.b_reg.out[14]$_DFFE_PP_  (.CLK(clknet_2_2__leaf_clk),
    .D(_092_),
    .QN(_027_));
 DFFHQNx1_ASAP7_75t_SL \dpath.b_reg.out[15]$_DFFE_PP_  (.CLK(clknet_2_2__leaf_clk),
    .D(_093_),
    .QN(_024_));
 DFFHQNx1_ASAP7_75t_SL \dpath.b_reg.out[1]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .D(_094_),
    .QN(_066_));
 DFFHQNx1_ASAP7_75t_SL \dpath.b_reg.out[2]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .D(_095_),
    .QN(_063_));
 DFFHQNx1_ASAP7_75t_SL \dpath.b_reg.out[3]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .D(_096_),
    .QN(_060_));
 DFFHQNx1_ASAP7_75t_SL \dpath.b_reg.out[4]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .D(_097_),
    .QN(_057_));
 DFFHQNx1_ASAP7_75t_SL \dpath.b_reg.out[5]$_DFFE_PP_  (.CLK(clknet_2_0__leaf_clk),
    .D(_098_),
    .QN(_054_));
 DFFHQNx1_ASAP7_75t_SL \dpath.b_reg.out[6]$_DFFE_PP_  (.CLK(clknet_2_0__leaf_clk),
    .D(_099_),
    .QN(_051_));
 DFFHQNx1_ASAP7_75t_SL \dpath.b_reg.out[7]$_DFFE_PP_  (.CLK(clknet_2_0__leaf_clk),
    .D(_100_),
    .QN(_048_));
 DFFHQNx1_ASAP7_75t_SL \dpath.b_reg.out[8]$_DFFE_PP_  (.CLK(clknet_2_0__leaf_clk),
    .D(_101_),
    .QN(_045_));
 DFFHQNx1_ASAP7_75t_SL \dpath.b_reg.out[9]$_DFFE_PP_  (.CLK(clknet_2_2__leaf_clk),
    .D(_102_),
    .QN(_042_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Left_52 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Left_53 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Left_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Left_55 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Left_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Left_57 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Left_58 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Left_59 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Left_60 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Left_61 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Left_62 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Left_63 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Left_64 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Left_65 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Left_66 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Left_67 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Left_68 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Left_69 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Left_70 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Left_71 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Left_72 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Left_73 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Left_74 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Left_75 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Left_76 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Left_77 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Left_78 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Left_79 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Left_80 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Left_81 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Left_82 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Left_83 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Left_84 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Left_85 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Left_86 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Left_87 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Left_88 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Left_89 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Left_90 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Left_91 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Left_92 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Left_93 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Left_94 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Left_95 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Left_96 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Left_97 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Left_98 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Left_99 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Left_100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Left_101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Left_102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Left_103 ();
 BUFx2_ASAP7_75t_L input16 (.A(req_msg[23]),
    .Y(net16));
 BUFx2_ASAP7_75t_L input17 (.A(req_msg[24]),
    .Y(net17));
 BUFx2_ASAP7_75t_L input18 (.A(req_msg[25]),
    .Y(net18));
 BUFx2_ASAP7_75t_L input19 (.A(req_msg[26]),
    .Y(net19));
 BUFx2_ASAP7_75t_L input20 (.A(req_msg[27]),
    .Y(net20));
 BUFx2_ASAP7_75t_L input21 (.A(req_msg[28]),
    .Y(net21));
 BUFx2_ASAP7_75t_L input22 (.A(req_msg[29]),
    .Y(net22));
 BUFx2_ASAP7_75t_L input23 (.A(req_msg[2]),
    .Y(net23));
 BUFx2_ASAP7_75t_L input24 (.A(req_msg[30]),
    .Y(net24));
 BUFx2_ASAP7_75t_L input25 (.A(req_msg[31]),
    .Y(net25));
 BUFx2_ASAP7_75t_L input26 (.A(req_msg[3]),
    .Y(net26));
 BUFx2_ASAP7_75t_L input27 (.A(req_msg[4]),
    .Y(net27));
 BUFx2_ASAP7_75t_L input28 (.A(req_msg[5]),
    .Y(net28));
 BUFx2_ASAP7_75t_L input29 (.A(req_msg[6]),
    .Y(net29));
 BUFx2_ASAP7_75t_L input30 (.A(req_msg[7]),
    .Y(net30));
 BUFx2_ASAP7_75t_L input31 (.A(req_msg[8]),
    .Y(net31));
 BUFx2_ASAP7_75t_L input32 (.A(req_msg[9]),
    .Y(net32));
 BUFx2_ASAP7_75t_L input33 (.A(req_val),
    .Y(net33));
 BUFx2_ASAP7_75t_L input34 (.A(reset),
    .Y(net34));
 BUFx2_ASAP7_75t_L input35 (.A(resp_rdy),
    .Y(net35));
 BUFx2_ASAP7_75t_L output36 (.A(net86),
    .Y(req_rdy));
 BUFx2_ASAP7_75t_L output37 (.A(net37),
    .Y(resp_msg[0]));
 BUFx2_ASAP7_75t_L output38 (.A(net38),
    .Y(resp_msg[10]));
 BUFx2_ASAP7_75t_L output39 (.A(net39),
    .Y(resp_msg[11]));
 BUFx2_ASAP7_75t_L output40 (.A(net40),
    .Y(resp_msg[12]));
 BUFx2_ASAP7_75t_L output41 (.A(net41),
    .Y(resp_msg[13]));
 BUFx2_ASAP7_75t_L output42 (.A(net42),
    .Y(resp_msg[14]));
 BUFx2_ASAP7_75t_L output43 (.A(net43),
    .Y(resp_msg[15]));
 BUFx2_ASAP7_75t_L output44 (.A(net44),
    .Y(resp_msg[1]));
 BUFx2_ASAP7_75t_L output45 (.A(net45),
    .Y(resp_msg[2]));
 BUFx2_ASAP7_75t_L output46 (.A(net46),
    .Y(resp_msg[3]));
 BUFx2_ASAP7_75t_L output47 (.A(net47),
    .Y(resp_msg[4]));
 BUFx2_ASAP7_75t_L output48 (.A(net48),
    .Y(resp_msg[5]));
 BUFx2_ASAP7_75t_L output49 (.A(net49),
    .Y(resp_msg[6]));
 BUFx2_ASAP7_75t_L output50 (.A(net50),
    .Y(resp_msg[7]));
 BUFx2_ASAP7_75t_L output51 (.A(net51),
    .Y(resp_msg[8]));
 BUFx2_ASAP7_75t_L output52 (.A(net52),
    .Y(resp_msg[9]));
 BUFx2_ASAP7_75t_L output53 (.A(net53),
    .Y(resp_val));
 BUFx6f_ASAP7_75t_L place83 (.A(_156_),
    .Y(net83));
 BUFx3_ASAP7_75t_L place82 (.A(_156_),
    .Y(net82));
 BUFx3_ASAP7_75t_L place84 (.A(_062_),
    .Y(net84));
 BUFx3_ASAP7_75t_L place85 (.A(_059_),
    .Y(net85));
 BUFx2_ASAP7_75t_R clkload2 (.A(clknet_2_3__leaf_clk));
 BUFx10_ASAP7_75t_SL clkload1 (.A(clknet_2_2__leaf_clk));
 BUFx2_ASAP7_75t_R clkload0 (.A(clknet_2_0__leaf_clk));
 BUFx4_ASAP7_75t_R clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Y(clknet_2_3__leaf_clk));
 BUFx4_ASAP7_75t_R clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Y(clknet_2_2__leaf_clk));
 BUFx4_ASAP7_75t_R clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Y(clknet_2_1__leaf_clk));
 BUFx3_ASAP7_75t_L place86 (.A(net36),
    .Y(net86));
 BUFx4_ASAP7_75t_R clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Y(clknet_2_0__leaf_clk));
 BUFx4_ASAP7_75t_R clkbuf_0_clk (.A(clk),
    .Y(clknet_0_clk));
endmodule
