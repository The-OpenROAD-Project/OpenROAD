module multi_sink (clk);
 input clk;

 DFF_X1 ff287 (.CK(clk));
 DFF_X1 ff286 (.CK(clk));
 DFF_X1 ff285 (.CK(clk));
 DFF_X1 ff284 (.CK(clk));
 DFF_X1 ff283 (.CK(clk));
 DFF_X1 ff282 (.CK(clk));
 DFF_X1 ff281 (.CK(clk));
 DFF_X1 ff280 (.CK(clk));
 DFF_X1 ff279 (.CK(clk));
 DFF_X1 ff278 (.CK(clk));
 DFF_X1 ff277 (.CK(clk));
 DFF_X1 ff276 (.CK(clk));
 DFF_X1 ff275 (.CK(clk));
 DFF_X1 ff274 (.CK(clk));
 DFF_X1 ff273 (.CK(clk));
 DFF_X1 ff272 (.CK(clk));
 DFF_X1 ff271 (.CK(clk));
 DFF_X1 ff270 (.CK(clk));
 DFF_X1 ff269 (.CK(clk));
 DFF_X1 ff268 (.CK(clk));
 DFF_X1 ff267 (.CK(clk));
 DFF_X1 ff266 (.CK(clk));
 DFF_X1 ff265 (.CK(clk));
 DFF_X1 ff264 (.CK(clk));
 DFF_X1 ff263 (.CK(clk));
 DFF_X1 ff262 (.CK(clk));
 DFF_X1 ff261 (.CK(clk));
 DFF_X1 ff260 (.CK(clk));
 DFF_X1 ff259 (.CK(clk));
 DFF_X1 ff258 (.CK(clk));
 DFF_X1 ff257 (.CK(clk));
 DFF_X1 ff256 (.CK(clk));
 DFF_X1 ff255 (.CK(clk));
 DFF_X1 ff254 (.CK(clk));
 DFF_X1 ff253 (.CK(clk));
 DFF_X1 ff252 (.CK(clk));
 DFF_X1 ff251 (.CK(clk));
 DFF_X1 ff250 (.CK(clk));
 DFF_X1 ff249 (.CK(clk));
 DFF_X1 ff248 (.CK(clk));
 DFF_X1 ff247 (.CK(clk));
 DFF_X1 ff246 (.CK(clk));
 DFF_X1 ff245 (.CK(clk));
 DFF_X1 ff244 (.CK(clk));
 DFF_X1 ff243 (.CK(clk));
 DFF_X1 ff242 (.CK(clk));
 DFF_X1 ff241 (.CK(clk));
 DFF_X1 ff240 (.CK(clk));
 DFF_X1 ff239 (.CK(clk));
 DFF_X1 ff238 (.CK(clk));
 DFF_X1 ff237 (.CK(clk));
 DFF_X1 ff236 (.CK(clk));
 DFF_X1 ff235 (.CK(clk));
 DFF_X1 ff234 (.CK(clk));
 DFF_X1 ff233 (.CK(clk));
 DFF_X1 ff232 (.CK(clk));
 DFF_X1 ff231 (.CK(clk));
 DFF_X1 ff230 (.CK(clk));
 DFF_X1 ff229 (.CK(clk));
 DFF_X1 ff228 (.CK(clk));
 DFF_X1 ff227 (.CK(clk));
 DFF_X1 ff226 (.CK(clk));
 DFF_X1 ff225 (.CK(clk));
 DFF_X1 ff224 (.CK(clk));
 DFF_X1 ff223 (.CK(clk));
 DFF_X1 ff222 (.CK(clk));
 DFF_X1 ff221 (.CK(clk));
 DFF_X1 ff220 (.CK(clk));
 DFF_X1 ff219 (.CK(clk));
 DFF_X1 ff218 (.CK(clk));
 DFF_X1 ff217 (.CK(clk));
 DFF_X1 ff216 (.CK(clk));
 DFF_X1 ff215 (.CK(clk));
 DFF_X1 ff214 (.CK(clk));
 DFF_X1 ff213 (.CK(clk));
 DFF_X1 ff212 (.CK(clk));
 DFF_X1 ff211 (.CK(clk));
 DFF_X1 ff210 (.CK(clk));
 DFF_X1 ff209 (.CK(clk));
 DFF_X1 ff208 (.CK(clk));
 DFF_X1 ff207 (.CK(clk));
 DFF_X1 ff206 (.CK(clk));
 DFF_X1 ff205 (.CK(clk));
 DFF_X1 ff204 (.CK(clk));
 DFF_X1 ff203 (.CK(clk));
 DFF_X1 ff202 (.CK(clk));
 DFF_X1 ff201 (.CK(clk));
 DFF_X1 ff200 (.CK(clk));
 DFF_X1 ff199 (.CK(clk));
 DFF_X1 ff198 (.CK(clk));
 DFF_X1 ff197 (.CK(clk));
 DFF_X1 ff196 (.CK(clk));
 DFF_X1 ff195 (.CK(clk));
 DFF_X1 ff194 (.CK(clk));
 DFF_X1 ff193 (.CK(clk));
 DFF_X1 ff192 (.CK(clk));
 DFF_X1 ff191 (.CK(clk));
 DFF_X1 ff190 (.CK(clk));
 DFF_X1 ff189 (.CK(clk));
 DFF_X1 ff188 (.CK(clk));
 DFF_X1 ff187 (.CK(clk));
 DFF_X1 ff186 (.CK(clk));
 DFF_X1 ff185 (.CK(clk));
 DFF_X1 ff184 (.CK(clk));
 DFF_X1 ff183 (.CK(clk));
 DFF_X1 ff182 (.CK(clk));
 DFF_X1 ff181 (.CK(clk));
 DFF_X1 ff180 (.CK(clk));
 DFF_X1 ff179 (.CK(clk));
 DFF_X1 ff178 (.CK(clk));
 DFF_X1 ff177 (.CK(clk));
 DFF_X1 ff176 (.CK(clk));
 DFF_X1 ff175 (.CK(clk));
 DFF_X1 ff174 (.CK(clk));
 DFF_X1 ff173 (.CK(clk));
 DFF_X1 ff172 (.CK(clk));
 DFF_X1 ff171 (.CK(clk));
 DFF_X1 ff170 (.CK(clk));
 DFF_X1 ff169 (.CK(clk));
 DFF_X1 ff168 (.CK(clk));
 DFF_X1 ff167 (.CK(clk));
 DFF_X1 ff166 (.CK(clk));
 DFF_X1 ff165 (.CK(clk));
 DFF_X1 ff164 (.CK(clk));
 DFF_X1 ff163 (.CK(clk));
 DFF_X1 ff162 (.CK(clk));
 DFF_X1 ff161 (.CK(clk));
 DFF_X1 ff160 (.CK(clk));
 DFF_X1 ff159 (.CK(clk));
 DFF_X1 ff158 (.CK(clk));
 DFF_X1 ff157 (.CK(clk));
 DFF_X1 ff156 (.CK(clk));
 DFF_X1 ff155 (.CK(clk));
 DFF_X1 ff154 (.CK(clk));
 DFF_X1 ff153 (.CK(clk));
 DFF_X1 ff152 (.CK(clk));
 DFF_X1 ff151 (.CK(clk));
 DFF_X1 ff150 (.CK(clk));
 DFF_X1 ff149 (.CK(clk));
 DFF_X1 ff148 (.CK(clk));
 DFF_X1 ff147 (.CK(clk));
 DFF_X1 ff146 (.CK(clk));
 DFF_X1 ff145 (.CK(clk));
 DFF_X1 ff144 (.CK(clk));
 DFF_X1 ff143 (.CK(clk));
 DFF_X1 ff142 (.CK(clk));
 DFF_X1 ff141 (.CK(clk));
 DFF_X1 ff140 (.CK(clk));
 DFF_X1 ff139 (.CK(clk));
 DFF_X1 ff138 (.CK(clk));
 DFF_X1 ff137 (.CK(clk));
 DFF_X1 ff136 (.CK(clk));
 DFF_X1 ff135 (.CK(clk));
 DFF_X1 ff134 (.CK(clk));
 DFF_X1 ff133 (.CK(clk));
 DFF_X1 ff132 (.CK(clk));
 DFF_X1 ff131 (.CK(clk));
 DFF_X1 ff130 (.CK(clk));
 DFF_X1 ff129 (.CK(clk));
 DFF_X1 ff125 (.CK(clk));
 DFF_X1 ff124 (.CK(clk));
 DFF_X1 ff123 (.CK(clk));
 DFF_X1 ff122 (.CK(clk));
 DFF_X1 ff121 (.CK(clk));
 DFF_X1 ff120 (.CK(clk));
 DFF_X1 ff119 (.CK(clk));
 DFF_X1 ff118 (.CK(clk));
 DFF_X1 ff117 (.CK(clk));
 DFF_X1 ff116 (.CK(clk));
 DFF_X1 ff115 (.CK(clk));
 DFF_X1 ff114 (.CK(clk));
 DFF_X1 ff113 (.CK(clk));
 DFF_X1 ff112 (.CK(clk));
 DFF_X1 ff111 (.CK(clk));
 DFF_X1 ff107 (.CK(clk));
 DFF_X1 ff106 (.CK(clk));
 DFF_X1 ff105 (.CK(clk));
 DFF_X1 ff104 (.CK(clk));
 DFF_X1 ff103 (.CK(clk));
 DFF_X1 ff102 (.CK(clk));
 DFF_X1 ff101 (.CK(clk));
 DFF_X1 ff100 (.CK(clk));
 DFF_X1 ff99 (.CK(clk));
 DFF_X1 ff98 (.CK(clk));
 DFF_X1 ff97 (.CK(clk));
 DFF_X1 ff96 (.CK(clk));
 DFF_X1 ff95 (.CK(clk));
 DFF_X1 ff94 (.CK(clk));
 DFF_X1 ff93 (.CK(clk));
 DFF_X1 ff92 (.CK(clk));
 DFF_X1 ff89 (.CK(clk));
 DFF_X1 ff88 (.CK(clk));
 DFF_X1 ff87 (.CK(clk));
 DFF_X1 ff86 (.CK(clk));
 DFF_X1 ff85 (.CK(clk));
 DFF_X1 ff84 (.CK(clk));
 DFF_X1 ff83 (.CK(clk));
 DFF_X1 ff82 (.CK(clk));
 DFF_X1 ff81 (.CK(clk));
 DFF_X1 ff80 (.CK(clk));
 DFF_X1 ff79 (.CK(clk));
 DFF_X1 ff78 (.CK(clk));
 DFF_X1 ff77 (.CK(clk));
 DFF_X1 ff76 (.CK(clk));
 DFF_X1 ff75 (.CK(clk));
 DFF_X1 ff74 (.CK(clk));
 DFF_X1 ff71 (.CK(clk));
 DFF_X1 ff70 (.CK(clk));
 DFF_X1 ff69 (.CK(clk));
 DFF_X1 ff68 (.CK(clk));
 DFF_X1 ff67 (.CK(clk));
 DFF_X1 ff66 (.CK(clk));
 DFF_X1 ff65 (.CK(clk));
 DFF_X1 ff64 (.CK(clk));
 DFF_X1 ff63 (.CK(clk));
 DFF_X1 ff62 (.CK(clk));
 DFF_X1 ff61 (.CK(clk));
 DFF_X1 ff60 (.CK(clk));
 DFF_X1 ff59 (.CK(clk));
 DFF_X1 ff58 (.CK(clk));
 DFF_X1 ff57 (.CK(clk));
 DFF_X1 ff56 (.CK(clk));
 DFF_X1 ff55 (.CK(clk));
 DFF_X1 ff54 (.CK(clk));
 DFF_X1 ff53 (.CK(clk));
 DFF_X1 ff52 (.CK(clk));
 DFF_X1 ff51 (.CK(clk));
 DFF_X1 ff50 (.CK(clk));
 DFF_X1 ff49 (.CK(clk));
 DFF_X1 ff48 (.CK(clk));
 DFF_X1 ff47 (.CK(clk));
 DFF_X1 ff46 (.CK(clk));
 DFF_X1 ff45 (.CK(clk));
 DFF_X1 ff44 (.CK(clk));
 DFF_X1 ff43 (.CK(clk));
 DFF_X1 ff42 (.CK(clk));
 DFF_X1 ff41 (.CK(clk));
 DFF_X1 ff40 (.CK(clk));
 DFF_X1 ff39 (.CK(clk));
 DFF_X1 ff38 (.CK(clk));
 DFF_X1 ff37 (.CK(clk));
 DFF_X1 ff36 (.CK(clk));
 DFF_X1 ff35 (.CK(clk));
 DFF_X1 ff34 (.CK(clk));
 DFF_X1 ff33 (.CK(clk));
 DFF_X1 ff32 (.CK(clk));
 DFF_X1 ff31 (.CK(clk));
 DFF_X1 ff30 (.CK(clk));
 DFF_X1 ff29 (.CK(clk));
 DFF_X1 ff28 (.CK(clk));
 DFF_X1 ff27 (.CK(clk));
 DFF_X1 ff26 (.CK(clk));
 DFF_X1 ff25 (.CK(clk));
 DFF_X1 ff24 (.CK(clk));
 DFF_X1 ff23 (.CK(clk));
 DFF_X1 ff22 (.CK(clk));
 DFF_X1 ff21 (.CK(clk));
 DFF_X1 ff20 (.CK(clk));
 DFF_X1 ff19 (.CK(clk));
 DFF_X1 ff18 (.CK(clk));
 DFF_X1 ff17 (.CK(clk));
 DFF_X1 ff16 (.CK(clk));
 DFF_X1 ff15 (.CK(clk));
 DFF_X1 ff14 (.CK(clk));
 DFF_X1 ff13 (.CK(clk));
 DFF_X1 ff12 (.CK(clk));
 DFF_X1 ff11 (.CK(clk));
 DFF_X1 ff10 (.CK(clk));
 DFF_X1 ff9 (.CK(clk));
 DFF_X1 ff8 (.CK(clk));
 DFF_X1 ff7 (.CK(clk));
 DFF_X1 ff6 (.CK(clk));
 DFF_X1 ff5 (.CK(clk));
 DFF_X1 ff4 (.CK(clk));

 hier_block h1(.childclk(clk));
   
 array_tile inst_0 (.clk(clk));
endmodule // multi_sink

module hier_block(childclk);
   input childclk;
 DFF_X1 ff3 (.CK(childclk));
 DFF_X1 ff2 (.CK(childclk));
 DFF_X1 ff1 (.CK(childclk));
 DFF_X1 ff0 (.CK(childclk));
endmodule // hier_block

