sky130_fd_sc_hs.tlef