../../../../test/sky130hd/sky130hd_std_cell.lef