module multi_sink (clk);
 input clk;

 wire gclk1;
 wire gclk3;
 wire gclk4;

 CLKGATE_X1 gclk1 (.CK(clk), .GCK(gclk1));
   DFF_X1 ff278 (.CK(gclk1));
   DFF_X1 ff277 (.CK(gclk1));
   DFF_X1 ff276 (.CK(gclk1));
   DFF_X1 ff275 (.CK(gclk1));
   DFF_X1 ff274 (.CK(gclk1));
   DFF_X1 ff273 (.CK(gclk1));
   DFF_X1 ff272 (.CK(gclk1));
   DFF_X1 ff271 (.CK(gclk1));
   DFF_X1 ff270 (.CK(gclk1));
   DFF_X1 ff260 (.CK(gclk1));
   DFF_X1 ff259 (.CK(gclk1));
   DFF_X1 ff258 (.CK(gclk1));
   DFF_X1 ff257 (.CK(gclk1));
   DFF_X1 ff256 (.CK(gclk1));
   DFF_X1 ff255 (.CK(gclk1));
   DFF_X1 ff254 (.CK(gclk1));
   DFF_X1 ff253 (.CK(gclk1));
   DFF_X1 ff252 (.CK(gclk1));
   DFF_X1 ff242 (.CK(gclk1));
   DFF_X1 ff241 (.CK(gclk1));
   DFF_X1 ff240 (.CK(gclk1));
   DFF_X1 ff239 (.CK(gclk1));
   DFF_X1 ff238 (.CK(gclk1));
   DFF_X1 ff237 (.CK(gclk1));
   DFF_X1 ff236 (.CK(gclk1));
   DFF_X1 ff235 (.CK(gclk1));
   DFF_X1 ff234 (.CK(gclk1));
   DFF_X1 ff224 (.CK(gclk1));
   DFF_X1 ff223 (.CK(gclk1));
   DFF_X1 ff222 (.CK(gclk1));
   DFF_X1 ff221 (.CK(gclk1));
   DFF_X1 ff220 (.CK(gclk1));
   DFF_X1 ff219 (.CK(gclk1));
   DFF_X1 ff218 (.CK(gclk1));
   DFF_X1 ff217 (.CK(gclk1));
   DFF_X1 ff216 (.CK(gclk1));
 CLKGATE_X1 gclk3 (.CK(gclk4), .GCK(gclk3));
 DFF_X1 ff287 (.CK(gclk3));
 DFF_X1 ff286 (.CK(gclk3));
 DFF_X1 ff285 (.CK(gclk3));
 DFF_X1 ff284 (.CK(gclk3));
 DFF_X1 ff283 (.CK(gclk3));
 DFF_X1 ff282 (.CK(gclk3));
 DFF_X1 ff281 (.CK(gclk3));
 DFF_X1 ff280 (.CK(gclk3));
 DFF_X1 ff279 (.CK(gclk3));
 DFF_X1 ff269 (.CK(gclk3));
 DFF_X1 ff268 (.CK(gclk3));
 DFF_X1 ff267 (.CK(gclk3));
 DFF_X1 ff266 (.CK(gclk3));
 DFF_X1 ff265 (.CK(gclk3));
 DFF_X1 ff264 (.CK(gclk3));
 DFF_X1 ff263 (.CK(gclk3));
 DFF_X1 ff262 (.CK(gclk3));
 DFF_X1 ff261 (.CK(gclk3));
 DFF_X1 ff251 (.CK(gclk3));
 DFF_X1 ff250 (.CK(gclk3));
 DFF_X1 ff249 (.CK(gclk3));
 DFF_X1 ff248 (.CK(gclk3));
 DFF_X1 ff247 (.CK(gclk3));
 DFF_X1 ff246 (.CK(gclk3));
 DFF_X1 ff245 (.CK(gclk3));
 DFF_X1 ff244 (.CK(gclk3));
 DFF_X1 ff243 (.CK(gclk3));
 DFF_X1 ff233 (.CK(gclk3));
 DFF_X1 ff232 (.CK(gclk3));
 DFF_X1 ff231 (.CK(gclk3));
 DFF_X1 ff230 (.CK(gclk3));
 DFF_X1 ff229 (.CK(gclk3));
 DFF_X1 ff228 (.CK(gclk3));
 DFF_X1 ff227 (.CK(gclk3));
 DFF_X1 ff226 (.CK(gclk3));
 DFF_X1 ff225 (.CK(gclk3));
 CLKGATE_X1 gclk4 (.CK(clk), .GCK(gclk4));
 DFF_X1 ff197 (.CK(gclk4));
 DFF_X1 ff196 (.CK(gclk4));
 DFF_X1 ff195 (.CK(gclk4));
 DFF_X1 ff194 (.CK(gclk4));
 DFF_X1 ff193 (.CK(gclk4));
 DFF_X1 ff192 (.CK(gclk4));
 DFF_X1 ff191 (.CK(gclk4));
 DFF_X1 ff190 (.CK(gclk4));
 DFF_X1 ff189 (.CK(gclk4));
 DFF_X1 ff179 (.CK(gclk4));
 DFF_X1 ff178 (.CK(gclk4));
 DFF_X1 ff177 (.CK(gclk4));
 DFF_X1 ff176 (.CK(gclk4));
 DFF_X1 ff175 (.CK(gclk4));
 DFF_X1 ff174 (.CK(gclk4));
 DFF_X1 ff173 (.CK(gclk4));
 DFF_X1 ff172 (.CK(gclk4));
 DFF_X1 ff171 (.CK(gclk4));
 DFF_X1 ff161 (.CK(gclk4));
 DFF_X1 ff160 (.CK(gclk4));
 DFF_X1 ff159 (.CK(gclk4));
 DFF_X1 ff158 (.CK(gclk4));
 DFF_X1 ff157 (.CK(gclk4));
 DFF_X1 ff156 (.CK(gclk4));
 DFF_X1 ff155 (.CK(gclk4));
 DFF_X1 ff154 (.CK(gclk4));
 DFF_X1 ff153 (.CK(gclk4));
 DFF_X1 ff215 (.CK(gclk4));
 DFF_X1 ff214 (.CK(gclk4));
 DFF_X1 ff213 (.CK(gclk4));
 DFF_X1 ff212 (.CK(gclk4));
 DFF_X1 ff211 (.CK(gclk4));
 DFF_X1 ff210 (.CK(gclk4));
 DFF_X1 ff209 (.CK(gclk4));
 DFF_X1 ff208 (.CK(gclk4));
 DFF_X1 ff207 (.CK(gclk4));

 hier_block h1(.childclk(clk));
endmodule // multi_sink

module hier_block(childclk);
   input childclk;

   wire gclk2;
   wire gclk5;

   CLKGATE_X1 gclk2 (.CK(childclk), .GCK(gclk2));
   DFF_X1 ff152 (.CK(gclk2));
   DFF_X1 ff151 (.CK(gclk2));
   DFF_X1 ff150 (.CK(gclk2));
   DFF_X1 ff149 (.CK(gclk2));
   DFF_X1 ff148 (.CK(gclk2));
   DFF_X1 ff147 (.CK(gclk2));
   DFF_X1 ff146 (.CK(gclk2));
   DFF_X1 ff145 (.CK(gclk2));
   DFF_X1 ff144 (.CK(gclk2));
   DFF_X1 ff170 (.CK(gclk2));
   DFF_X1 ff169 (.CK(gclk2));
   DFF_X1 ff168 (.CK(gclk2));
   DFF_X1 ff167 (.CK(gclk2));
   DFF_X1 ff166 (.CK(gclk2));
   DFF_X1 ff165 (.CK(gclk2));
   DFF_X1 ff164 (.CK(gclk2));
   DFF_X1 ff163 (.CK(gclk2));
   DFF_X1 ff162 (.CK(gclk2));
   DFF_X1 ff188 (.CK(gclk2));
   DFF_X1 ff187 (.CK(gclk2));
   DFF_X1 ff186 (.CK(gclk2));
   DFF_X1 ff185 (.CK(gclk2));
   DFF_X1 ff184 (.CK(gclk2));
   DFF_X1 ff183 (.CK(gclk2));
   DFF_X1 ff182 (.CK(gclk2));
   DFF_X1 ff181 (.CK(gclk2));
   DFF_X1 ff180 (.CK(gclk2));
   DFF_X1 ff206 (.CK(gclk2));
   DFF_X1 ff205 (.CK(gclk2));
   DFF_X1 ff204 (.CK(gclk2));
   DFF_X1 ff203 (.CK(gclk2));
   DFF_X1 ff202 (.CK(gclk2));
   DFF_X1 ff201 (.CK(gclk2));
   DFF_X1 ff200 (.CK(gclk2));
   DFF_X1 ff199 (.CK(gclk2));
   DFF_X1 ff198 (.CK(gclk2));
   CLKGATE_X1 gclk5 (.CK(childclk), .GCK(gclk5));
   DFF_X1 ff143 (.CK(gclk5));
   DFF_X1 ff142 (.CK(gclk5));
   DFF_X1 ff141 (.CK(gclk5));
   DFF_X1 ff140 (.CK(gclk5));
   DFF_X1 ff139 (.CK(gclk5));
   DFF_X1 ff138 (.CK(gclk5));
   DFF_X1 ff137 (.CK(gclk5));
   DFF_X1 ff136 (.CK(gclk5));
   DFF_X1 ff135 (.CK(gclk5));
   DFF_X1 ff134 (.CK(gclk5));
   DFF_X1 ff133 (.CK(gclk5));
   DFF_X1 ff132 (.CK(gclk5));
   DFF_X1 ff131 (.CK(gclk5));
   DFF_X1 ff130 (.CK(gclk5));
   DFF_X1 ff129 (.CK(gclk5));
   DFF_X1 ff125 (.CK(gclk5));
   DFF_X1 ff124 (.CK(gclk5));
   DFF_X1 ff123 (.CK(gclk5));
   DFF_X1 ff122 (.CK(gclk5));
   DFF_X1 ff121 (.CK(gclk5));
   DFF_X1 ff120 (.CK(gclk5));
   DFF_X1 ff119 (.CK(gclk5));
   DFF_X1 ff118 (.CK(gclk5));
   DFF_X1 ff117 (.CK(gclk5));
   DFF_X1 ff116 (.CK(gclk5));
   DFF_X1 ff115 (.CK(gclk5));
   DFF_X1 ff114 (.CK(gclk5));
   DFF_X1 ff113 (.CK(gclk5));
   DFF_X1 ff112 (.CK(gclk5));
   DFF_X1 ff111 (.CK(gclk5));
   DFF_X1 ff107 (.CK(gclk5));
   DFF_X1 ff106 (.CK(gclk5));
   DFF_X1 ff105 (.CK(gclk5));
   DFF_X1 ff104 (.CK(gclk5));
   DFF_X1 ff103 (.CK(gclk5));
   DFF_X1 ff102 (.CK(gclk5));
   DFF_X1 ff101 (.CK(gclk5));
   DFF_X1 ff100 (.CK(gclk5));
   DFF_X1 ff99 (.CK(gclk5));
   DFF_X1 ff98 (.CK(gclk5));
   DFF_X1 ff97 (.CK(gclk5));
   DFF_X1 ff96 (.CK(gclk5));
   DFF_X1 ff95 (.CK(gclk5));
   DFF_X1 ff94 (.CK(gclk5));
   DFF_X1 ff93 (.CK(gclk5));
   DFF_X1 ff92 (.CK(gclk5));
   DFF_X1 ff89 (.CK(gclk5));
   DFF_X1 ff88 (.CK(gclk5));
   DFF_X1 ff87 (.CK(gclk5));
   DFF_X1 ff86 (.CK(gclk5));
   DFF_X1 ff85 (.CK(gclk5));
   DFF_X1 ff84 (.CK(gclk5));
   DFF_X1 ff83 (.CK(gclk5));
   DFF_X1 ff82 (.CK(gclk5));
   DFF_X1 ff81 (.CK(gclk5));
   DFF_X1 ff80 (.CK(gclk5));
   DFF_X1 ff79 (.CK(gclk5));
   DFF_X1 ff78 (.CK(gclk5));
   DFF_X1 ff77 (.CK(gclk5));
   DFF_X1 ff76 (.CK(gclk5));
   DFF_X1 ff75 (.CK(gclk5));
   DFF_X1 ff74 (.CK(gclk5));
   DFF_X1 ff71 (.CK(gclk5));
   DFF_X1 ff70 (.CK(gclk5));
   DFF_X1 ff69 (.CK(gclk5));
   DFF_X1 ff68 (.CK(gclk5));
   DFF_X1 ff67 (.CK(gclk5));
   DFF_X1 ff66 (.CK(gclk5));
   DFF_X1 ff65 (.CK(gclk5));
   DFF_X1 ff64 (.CK(gclk5));
   DFF_X1 ff63 (.CK(gclk5));
   DFF_X1 ff62 (.CK(gclk5));
   DFF_X1 ff61 (.CK(gclk5));
   DFF_X1 ff60 (.CK(gclk5));
   DFF_X1 ff59 (.CK(gclk5));
   DFF_X1 ff58 (.CK(gclk5));
   DFF_X1 ff57 (.CK(gclk5));
   DFF_X1 ff56 (.CK(gclk5));
   DFF_X1 ff55 (.CK(gclk5));
   DFF_X1 ff54 (.CK(gclk5));
   DFF_X1 ff53 (.CK(gclk5));
   DFF_X1 ff52 (.CK(gclk5));
   DFF_X1 ff51 (.CK(gclk5));
   DFF_X1 ff50 (.CK(gclk5));
   DFF_X1 ff49 (.CK(gclk5));
   DFF_X1 ff48 (.CK(gclk5));
   DFF_X1 ff47 (.CK(gclk5));
   DFF_X1 ff46 (.CK(gclk5));
   DFF_X1 ff45 (.CK(gclk5));
   DFF_X1 ff44 (.CK(gclk5));
   DFF_X1 ff43 (.CK(gclk5));
   DFF_X1 ff42 (.CK(gclk5));
   DFF_X1 ff41 (.CK(gclk5));
   DFF_X1 ff40 (.CK(gclk5));
   DFF_X1 ff39 (.CK(gclk5));
   DFF_X1 ff38 (.CK(gclk5));
   DFF_X1 ff37 (.CK(gclk5));
   DFF_X1 ff36 (.CK(gclk5));
   DFF_X1 ff35 (.CK(gclk5));
   DFF_X1 ff34 (.CK(gclk5));
   DFF_X1 ff33 (.CK(gclk5));
   DFF_X1 ff32 (.CK(gclk5));
   DFF_X1 ff31 (.CK(gclk5));
   DFF_X1 ff30 (.CK(gclk5));
   DFF_X1 ff29 (.CK(gclk5));
   DFF_X1 ff28 (.CK(gclk5));
   DFF_X1 ff27 (.CK(gclk5));
   DFF_X1 ff26 (.CK(gclk5));
   DFF_X1 ff25 (.CK(gclk5));
   DFF_X1 ff24 (.CK(gclk5));
   DFF_X1 ff23 (.CK(gclk5));
   DFF_X1 ff22 (.CK(gclk5));
   DFF_X1 ff21 (.CK(gclk5));
   DFF_X1 ff20 (.CK(gclk5));
   DFF_X1 ff19 (.CK(gclk5));
   DFF_X1 ff18 (.CK(gclk5));
   DFF_X1 ff17 (.CK(gclk5));
   DFF_X1 ff16 (.CK(gclk5));
   DFF_X1 ff15 (.CK(gclk5));
   DFF_X1 ff14 (.CK(gclk5));
   DFF_X1 ff13 (.CK(gclk5));
   DFF_X1 ff12 (.CK(gclk5));
   DFF_X1 ff11 (.CK(gclk5));
   DFF_X1 ff10 (.CK(gclk5));
   DFF_X1 ff9 (.CK(gclk5));
   DFF_X1 ff8 (.CK(gclk5));
   DFF_X1 ff7 (.CK(gclk5));
   DFF_X1 ff6 (.CK(gclk5));
   DFF_X1 ff5 (.CK(gclk5));
   DFF_X1 ff4 (.CK(gclk5));
   DFF_X1 ff3 (.CK(gclk5));
   DFF_X1 ff2 (.CK(gclk5));
   DFF_X1 ff1 (.CK(gclk5));
   DFF_X1 \ff0/name (.CK(gclk5));
 
endmodule // hier_block1

