VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

SITE DoubleHeightSite
  SYMMETRY X Y ;
  CLASS core ;
  SIZE 0.19 BY 2.8 ;
END DoubleHeightSite


SITE TripleHeightSite
  SYMMETRY Y ;
  CLASS core ;
  SIZE 0.19 BY 4.2 ;
END TripleHeightSite

MACRO MOCK_SINGLE
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2_X1 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT VERTICAL_EDGE_1 ;
    EDGETYPE RIGHT VERTICAL_EDGE_1 ; " ;
  PIN A1 
  END A1
  PIN A2 
  END A2
  PIN ZN 
  END ZN
  PIN VDD 
  END VDD
  PIN VSS 
  END VSS
END MOCK_SINGLE

MACRO MOCK_DOUBLE
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2_X1 0 0 ;
  SIZE 0.76 BY 2.8 ;
  SYMMETRY X Y ;
  SITE DoubleHeightSite ;
  PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT VERTICAL_EDGE_1 CELLROW 1 ;
    EDGETYPE LEFT VERTICAL_EDGE_2 CELLROW 2 ;
    EDGETYPE RIGHT VERTICAL_EDGE_1 CELLROW 1 ;
    EDGETYPE RIGHT VERTICAL_EDGE_2 CELLROW 2 ; " ;
  PIN A1 
  END A1
  PIN A2 
  END A2
  PIN ZN 
  END ZN
  PIN VDD 
  END VDD
  PIN VSS 
  END VSS
END MOCK_DOUBLE

MACRO MOCK_TRIPLE
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2_X1 0 0 ;
  SIZE 0.76 BY 4.2 ;
  SYMMETRY X Y ;
  SITE TripleHeightSite ;
  PIN A1 
  END A1
  PIN A2 
  END A2
  PIN ZN 
  END ZN
  PIN VDD 
  END VDD
  PIN VSS 
  END VSS
END MOCK_TRIPLE
