sky130_fd_sc_hd_merged.lef