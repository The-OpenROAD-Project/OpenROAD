VERSION	5.7 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  LAYER contactResistance REAL ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MANUFACTURINGGRID 0.0025 ;
LAYER poly
  TYPE MASTERSLICE ;
END poly

LAYER contact
  TYPE CUT ;
  SPACING 0.075 ;
  PROPERTY contactResistance 10.5 ;
END contact

LAYER metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.19 ;
  WIDTH 0.065 ;
  SPACING 0.065 ;
  RESISTANCE RPERSQ 0.38 ;
END metal1

LAYER via1
  TYPE CUT ;
  SPACING 0.075 ;
  PROPERTY contactResistance 5.69 ;
END via1

LAYER metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.19 ;
  WIDTH 0.07 ;
  SPACING 0.075 ;
  RESISTANCE RPERSQ 0.25 ;
END metal2

LAYER via2
  TYPE CUT ;
  SPACING 0.085 ;
  PROPERTY contactResistance 11.39 ;
END via2

LAYER metal3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.19 ;
  WIDTH 0.07 ;
  SPACING 0.07 ;
  RESISTANCE RPERSQ 0.25 ;
END metal3

LAYER via3
  TYPE CUT ;
  SPACING 0.085 ;
  PROPERTY contactResistance 16.73 ;
END via3

LAYER metal4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.285 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  RESISTANCE RPERSQ 0.25 ;
END metal4

LAYER via4
  TYPE CUT ;
  SPACING 0.16 ;
  PROPERTY contactResistance 21.44 ;
END via4

LAYER metal5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.285 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  RESISTANCE RPERSQ 0.25 ;
END metal5

LAYER via5
  TYPE CUT ;
  SPACING 0.16 ;
  PROPERTY contactResistance 24.08 ;
END via5

LAYER metal6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.285 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  RESISTANCE RPERSQ 0.25 ;
END metal6

LAYER via6
  TYPE CUT ;
  SPACING 0.16 ;
  PROPERTY contactResistance 11.39 ;
END via6

LAYER metal7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.855 ;
  WIDTH 0.4 ;
  SPACING 0.4 ;
  RESISTANCE RPERSQ 0.25 ;
END metal7

LAYER via7
  TYPE CUT ;
  SPACING 0.44 ;
  PROPERTY contactResistance 5.69 ;
END via7

LAYER metal8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.855 ;
  WIDTH 0.4 ;
  SPACING 0.4 ;
  RESISTANCE RPERSQ 0.25 ;
END metal8

LAYER via8
  TYPE CUT ;
  SPACING 0.44 ;
  PROPERTY contactResistance 16.73 ;
END via8

LAYER metal9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1.71 ;
  WIDTH 0.8 ;
  SPACING 0.8 ;
  RESISTANCE RPERSQ 0.21 ;
END metal9

LAYER via9
  TYPE CUT ;
  SPACING 0.88 ;
  PROPERTY contactResistance 21.44 ;
END via9

LAYER metal10
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 1.71 ;
  WIDTH 0.8 ;
  SPACING 0.8 ;
  RESISTANCE RPERSQ 0.21 ;
END metal10

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA M2_M1_via DEFAULT
  LAYER metal1 ;
    RECT -0.0675 -0.0325 0.0675 0.0325 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal2 ;
    RECT -0.035 -0.0675 0.035 0.0675 ;
END M2_M1_via

VIA M3_M2_via DEFAULT
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END M3_M2_via

VIA M4_M3_via DEFAULT
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M4_M3_via

VIA M5_M4_via DEFAULT
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M5_M4_via

VIA M6_M5_via DEFAULT
  LAYER metal5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M6_M5_via

VIA M7_M6_via DEFAULT
  LAYER metal6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END M7_M6_via

VIA M8_M7_via DEFAULT
  LAYER metal7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END M8_M7_via

VIA M9_M8_via DEFAULT
  LAYER metal8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END M9_M8_via

VIA M10_M9_via DEFAULT
  LAYER metal9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER metal10 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END M10_M9_via

VIA M2_M1_viaB DEFAULT
  LAYER metal1 ;
    RECT -0.0675 -0.0325 0.0675 0.0325 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal2 ;
    RECT -0.0675 -0.035 0.0675 0.035 ;
END M2_M1_viaB

VIA M2_M1_viaC DEFAULT
  LAYER metal1 ;
    RECT -0.0325 -0.0675 0.0325 0.0675 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal2 ;
    RECT -0.035 -0.0675 0.035 0.0675 ;
END M2_M1_viaC

VIA M3_M2_viaB DEFAULT
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END M3_M2_viaB

VIA M3_M2_viaC DEFAULT
  LAYER metal2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END M3_M2_viaC

VIA M4_M3_viaB DEFAULT
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M4_M3_viaB

VIARULE M2_M1 GENERATE
  LAYER metal1 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal2 ;
    ENCLOSURE 0 0.035 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
    SPACING 0.14 BY 0.14 ;
END M2_M1

VIARULE M3_M2 GENERATE
  LAYER metal2 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.155 BY 0.155 ;
END M3_M2

VIARULE M4_M3 GENERATE
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal4 ;
    ENCLOSURE 0 0 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.155 BY 0.155 ;
END M4_M3

VIARULE M5_M4 GENERATE
  LAYER metal4 ;
    ENCLOSURE 0 0 ;
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END M5_M4

VIARULE M6_M5 GENERATE
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END M6_M5

VIARULE M7_M6 GENERATE
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
  LAYER metal7 ;
    ENCLOSURE 0.13 0.13 ;
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END M7_M6

VIARULE M8_M7 GENERATE
  LAYER metal7 ;
    ENCLOSURE 0 0 ;
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.84 BY 0.84 ;
END M8_M7

VIARULE M9_M8 GENERATE
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
  LAYER metal9 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.84 BY 0.84 ;
END M9_M8

VIARULE M10_M9 GENERATE
  LAYER metal9 ;
    ENCLOSURE 0 0 ;
  LAYER metal10 ;
    ENCLOSURE 0 0 ;
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
    SPACING 1.68 BY 1.68 ;
END M10_M9

VIARULE M1_POLY GENERATE
  LAYER poly ;
    ENCLOSURE 0 0 ;
  LAYER metal1 ;
    ENCLOSURE 0 0.035 ;
  LAYER contact ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
    SPACING 0.14 BY 0.14 ;
END M1_POLY

SPACING
  SAMENET metal1 metal1 0.065 ;
  SAMENET metal2 metal2 0.07 ;
  SAMENET metal6 metal6 0.14 ;
  SAMENET metal5 metal5 0.14 ;
  SAMENET metal4 metal4 0.14 ;
  SAMENET metal3 metal3 0.07 ;
  SAMENET metal7 metal7 0.4 ;
  SAMENET metal8 metal8 0.4 ;
  SAMENET metal9 metal9 0.8 ;
  SAMENET metal10 metal10 0.8 ;
END SPACING

SITE CoreSite
  CLASS CORE ;
  SIZE 0.38 BY 1.71 ;
END CoreSite

MACRO in01s01
    CLASS CORE ;
    FOREIGN in01s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.695 0.150 0.825 1.255 ;
        RECT 0.625 0.150 0.885 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.315 0.340 0.51 0.405 ;
        END
    END a
END in01s01

MACRO in01s02
    CLASS CORE ;
    FOREIGN in01s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.280 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.150 1.65 1.255 ;
        RECT 1.250 0.150 1.77 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.340 1.02 0.405 ;
        END
    END a
END in01s02

MACRO in01s03
    CLASS CORE ;
    FOREIGN in01s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.150 1.945 1.255 ;
        RECT 1.460 0.150 2.11 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.340 1.19 0.405 ;
        END
    END a
END in01s03

MACRO in01s04
    CLASS CORE ;
    FOREIGN in01s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.040 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.150 2.18 1.255 ;
        RECT 1.665 0.150 2.38 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.840 0.340 1.36 0.405 ;
        END
    END a
END in01s04

MACRO in01s06
    CLASS CORE ;
    FOREIGN in01s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.150 2.475 1.255 ;
        RECT 1.875 0.150 2.655 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.945 0.340 1.53 0.405 ;
        END
    END a
END in01s06

MACRO in01s08
    CLASS CORE ;
    FOREIGN in01s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.315 0.150 2.77 1.255 ;
        RECT 2.085 0.150 2.995 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.050 0.340 1.7 0.405 ;
        END
    END a
END in01s08

MACRO in01s10
    CLASS CORE ;
    FOREIGN in01s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.180 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.550 0.150 3.005 1.255 ;
        RECT 2.290 0.150 3.265 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.155 0.340 1.87 0.405 ;
        END
    END a
END in01s10

MACRO in01s20
    CLASS CORE ;
    FOREIGN in01s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.245 0.150 3.83 1.255 ;
        RECT 2.915 0.150 4.15 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.470 0.340 2.38 0.405 ;
        END
    END a
END in01s20

MACRO in01s40
    CLASS CORE ;
    FOREIGN in01s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.220 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.400 0.150 5.245 1.255 ;
        RECT 3.960 0.150 5.65 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.995 0.340 3.23 0.405 ;
        END
    END a
END in01s40

MACRO in01s80
    CLASS CORE ;
    FOREIGN in01s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.880 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.025 0.150 7.13 1.255 ;
        RECT 5.415 0.150 7.755 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.730 0.340 4.485 0.405 ;
        END
    END a
END in01s80

MACRO in01m01
    CLASS CORE ;
    FOREIGN in01m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.695 0.150 0.825 1.255 ;
        RECT 0.625 0.150 0.885 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.315 0.340 0.51 0.405 ;
        END
    END a
END in01m01

MACRO in01m02
    CLASS CORE ;
    FOREIGN in01m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.280 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.150 1.65 1.255 ;
        RECT 1.250 0.150 1.77 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.340 1.02 0.405 ;
        END
    END a
END in01m02

MACRO in01m03
    CLASS CORE ;
    FOREIGN in01m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.150 1.945 1.255 ;
        RECT 1.460 0.150 2.11 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.340 1.19 0.405 ;
        END
    END a
END in01m03

MACRO in01m04
    CLASS CORE ;
    FOREIGN in01m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.040 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.150 2.18 1.255 ;
        RECT 1.665 0.150 2.38 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.840 0.340 1.36 0.405 ;
        END
    END a
END in01m04

MACRO in01m06
    CLASS CORE ;
    FOREIGN in01m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.150 2.475 1.255 ;
        RECT 1.875 0.150 2.655 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.945 0.340 1.53 0.405 ;
        END
    END a
END in01m06

MACRO in01m08
    CLASS CORE ;
    FOREIGN in01m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.315 0.150 2.77 1.255 ;
        RECT 2.085 0.150 2.995 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.050 0.340 1.7 0.405 ;
        END
    END a
END in01m08

MACRO in01m10
    CLASS CORE ;
    FOREIGN in01m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.180 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.550 0.150 3.005 1.255 ;
        RECT 2.290 0.150 3.265 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.155 0.340 1.87 0.405 ;
        END
    END a
END in01m10

MACRO in01m20
    CLASS CORE ;
    FOREIGN in01m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.245 0.150 3.83 1.255 ;
        RECT 2.915 0.150 4.15 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.470 0.340 2.38 0.405 ;
        END
    END a
END in01m20

MACRO in01m40
    CLASS CORE ;
    FOREIGN in01m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.220 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.400 0.150 5.245 1.255 ;
        RECT 3.960 0.150 5.65 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.995 0.340 3.23 0.405 ;
        END
    END a
END in01m40

MACRO in01m80
    CLASS CORE ;
    FOREIGN in01m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.880 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.025 0.150 7.13 1.255 ;
        RECT 5.415 0.150 7.755 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.730 0.340 4.485 0.405 ;
        END
    END a
END in01m80

MACRO in01f01
    CLASS CORE ;
    FOREIGN in01f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.695 0.150 0.825 1.255 ;
        RECT 0.625 0.150 0.885 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.315 0.340 0.51 0.405 ;
        END
    END a
END in01f01

MACRO in01f02
    CLASS CORE ;
    FOREIGN in01f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.280 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.150 1.65 1.255 ;
        RECT 1.250 0.150 1.77 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.340 1.02 0.405 ;
        END
    END a
END in01f02

MACRO in01f03
    CLASS CORE ;
    FOREIGN in01f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.150 1.945 1.255 ;
        RECT 1.460 0.150 2.11 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.340 1.19 0.405 ;
        END
    END a
END in01f03

MACRO in01f04
    CLASS CORE ;
    FOREIGN in01f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.040 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.150 2.18 1.255 ;
        RECT 1.665 0.150 2.38 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.840 0.340 1.36 0.405 ;
        END
    END a
END in01f04

MACRO in01f06
    CLASS CORE ;
    FOREIGN in01f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.150 2.475 1.255 ;
        RECT 1.875 0.150 2.655 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.945 0.340 1.53 0.405 ;
        END
    END a
END in01f06

MACRO in01f08
    CLASS CORE ;
    FOREIGN in01f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.315 0.150 2.77 1.255 ;
        RECT 2.085 0.150 2.995 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.050 0.340 1.7 0.405 ;
        END
    END a
END in01f08

MACRO in01f10
    CLASS CORE ;
    FOREIGN in01f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.180 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.550 0.150 3.005 1.255 ;
        RECT 2.290 0.150 3.265 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.155 0.340 1.87 0.405 ;
        END
    END a
END in01f10

MACRO in01f20
    CLASS CORE ;
    FOREIGN in01f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.245 0.150 3.83 1.255 ;
        RECT 2.915 0.150 4.15 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.470 0.340 2.38 0.405 ;
        END
    END a
END in01f20

MACRO in01f40
    CLASS CORE ;
    FOREIGN in01f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.220 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.400 0.150 5.245 1.255 ;
        RECT 3.960 0.150 5.65 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.995 0.340 3.23 0.405 ;
        END
    END a
END in01f40

MACRO in01f80
    CLASS CORE ;
    FOREIGN in01f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.880 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.025 0.150 7.13 1.255 ;
        RECT 5.415 0.150 7.755 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.730 0.340 4.485 0.405 ;
        END
    END a
END in01f80

MACRO na02s01
    CLASS CORE ;
    FOREIGN na02s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.450 0.110 0.58 1.215 ;
        RECT 0.430 0.725 0.625 1.245 ;
        RECT 0.450 0.110 0.905 0.175 ;
        RECT 0.805 0.110 0.935 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.070 0.535 0.33 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.645 0.540 0.905 0.67 ;
        END
    END b
END na02s01

MACRO na02s02
    CLASS CORE ;
    FOREIGN na02s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.800 0.110 2.19 1.215 ;
        RECT 1.710 0.725 2.49 1.245 ;
        RECT 1.800 0.110 3.62 0.175 ;
        RECT 3.210 0.110 3.6 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.270 0.535 1.44 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.540 3.62 0.67 ;
        END
    END b
END na02s02

MACRO na02s03
    CLASS CORE ;
    FOREIGN na02s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.250 0.110 2.77 1.215 ;
        RECT 2.140 0.725 3.18 1.245 ;
        RECT 2.250 0.110 4.525 0.175 ;
        RECT 4.015 0.110 4.535 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.340 0.535 1.77 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.225 0.540 4.525 0.67 ;
        END
    END b
END na02s03

MACRO na02s04
    CLASS CORE ;
    FOREIGN na02s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.840 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.700 0.110 3.285 1.215 ;
        RECT 2.565 0.725 3.8 1.245 ;
        RECT 2.700 0.110 5.43 0.175 ;
        RECT 4.815 0.110 5.4 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.405 0.535 2.095 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.870 0.540 5.43 0.67 ;
        END
    END b
END na02s04

MACRO na02s06
    CLASS CORE ;
    FOREIGN na02s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.300 0.110 4.015 1.215 ;
        RECT 3.135 0.725 4.63 1.245 ;
        RECT 3.300 0.110 6.615 0.175 ;
        RECT 5.885 0.110 6.6 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.495 0.535 2.575 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.730 0.540 6.615 0.67 ;
        END
    END b
END na02s06

MACRO na02s08
    CLASS CORE ;
    FOREIGN na02s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.880 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.900 0.110 4.745 1.215 ;
        RECT 3.705 0.725 5.46 1.245 ;
        RECT 3.900 0.110 7.8 0.175 ;
        RECT 6.955 0.110 7.8 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.585 0.535 3.055 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.590 0.540 7.865 0.67 ;
        END
    END b
END na02s08

MACRO na02s10
    CLASS CORE ;
    FOREIGN na02s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.020 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.350 0.110 5.325 1.215 ;
        RECT 4.135 0.725 6.085 1.245 ;
        RECT 4.350 0.110 8.705 0.175 ;
        RECT 7.760 0.110 8.735 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.655 0.535 3.385 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.235 0.540 8.705 0.67 ;
        END
    END b
END na02s10

MACRO na02s20
    CLASS CORE ;
    FOREIGN na02s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.150 0.110 7.515 1.215 ;
        RECT 5.845 0.725 8.64 1.245 ;
        RECT 6.150 0.110 12.325 0.175 ;
        RECT 10.970 0.110 12.335 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.535 4.825 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.815 0.540 12.325 0.67 ;
        END
    END b
END na02s20

MACRO na02s40
    CLASS CORE ;
    FOREIGN na02s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.550 0.110 10.435 1.215 ;
        RECT 8.125 0.725 11.96 1.245 ;
        RECT 8.550 0.110 17.13 0.175 ;
        RECT 15.250 0.110 17.135 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.285 0.535 6.68 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.255 0.540 17.195 0.67 ;
        END
    END b
END na02s40

MACRO na02s80
    CLASS CORE ;
    FOREIGN na02s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.400 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.000 0.110 14.6 1.215 ;
        RECT 11.400 0.725 16.795 1.245 ;
        RECT 12.000 0.110 24.025 0.175 ;
        RECT 21.400 0.110 24.0 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.800 0.535 9.405 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 17.200 0.540 24.09 0.67 ;
        END
    END b
END na02s80

MACRO na02m01
    CLASS CORE ;
    FOREIGN na02m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.450 0.110 0.58 1.215 ;
        RECT 0.430 0.725 0.625 1.245 ;
        RECT 0.450 0.110 0.905 0.175 ;
        RECT 0.805 0.110 0.935 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.070 0.535 0.33 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.645 0.540 0.905 0.67 ;
        END
    END b
END na02m01

MACRO na02m02
    CLASS CORE ;
    FOREIGN na02m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.800 0.110 2.19 1.215 ;
        RECT 1.710 0.725 2.49 1.245 ;
        RECT 1.800 0.110 3.62 0.175 ;
        RECT 3.210 0.110 3.6 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.270 0.535 1.44 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.540 3.62 0.67 ;
        END
    END b
END na02m02

MACRO na02m03
    CLASS CORE ;
    FOREIGN na02m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.250 0.110 2.77 1.215 ;
        RECT 2.140 0.725 3.18 1.245 ;
        RECT 2.250 0.110 4.525 0.175 ;
        RECT 4.015 0.110 4.535 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.340 0.535 1.77 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.225 0.540 4.525 0.67 ;
        END
    END b
END na02m03

MACRO na02m04
    CLASS CORE ;
    FOREIGN na02m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.840 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.700 0.110 3.285 1.215 ;
        RECT 2.565 0.725 3.8 1.245 ;
        RECT 2.700 0.110 5.43 0.175 ;
        RECT 4.815 0.110 5.4 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.405 0.535 2.095 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.870 0.540 5.43 0.67 ;
        END
    END b
END na02m04

MACRO na02m06
    CLASS CORE ;
    FOREIGN na02m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.300 0.110 4.015 1.215 ;
        RECT 3.135 0.725 4.63 1.245 ;
        RECT 3.300 0.110 6.615 0.175 ;
        RECT 5.885 0.110 6.6 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.495 0.535 2.575 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.730 0.540 6.615 0.67 ;
        END
    END b
END na02m06

MACRO na02m08
    CLASS CORE ;
    FOREIGN na02m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.880 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.900 0.110 4.745 1.215 ;
        RECT 3.705 0.725 5.46 1.245 ;
        RECT 3.900 0.110 7.8 0.175 ;
        RECT 6.955 0.110 7.8 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.585 0.535 3.055 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.590 0.540 7.865 0.67 ;
        END
    END b
END na02m08

MACRO na02m10
    CLASS CORE ;
    FOREIGN na02m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.020 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.350 0.110 5.325 1.215 ;
        RECT 4.135 0.725 6.085 1.245 ;
        RECT 4.350 0.110 8.705 0.175 ;
        RECT 7.760 0.110 8.735 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.655 0.535 3.385 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.235 0.540 8.705 0.67 ;
        END
    END b
END na02m10

MACRO na02m20
    CLASS CORE ;
    FOREIGN na02m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.150 0.110 7.515 1.215 ;
        RECT 5.845 0.725 8.64 1.245 ;
        RECT 6.150 0.110 12.325 0.175 ;
        RECT 10.970 0.110 12.335 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.535 4.825 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.815 0.540 12.325 0.67 ;
        END
    END b
END na02m20

MACRO na02m40
    CLASS CORE ;
    FOREIGN na02m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.550 0.110 10.435 1.215 ;
        RECT 8.125 0.725 11.96 1.245 ;
        RECT 8.550 0.110 17.13 0.175 ;
        RECT 15.250 0.110 17.135 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.285 0.535 6.68 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.255 0.540 17.195 0.67 ;
        END
    END b
END na02m40

MACRO na02m80
    CLASS CORE ;
    FOREIGN na02m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.400 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.000 0.110 14.6 1.215 ;
        RECT 11.400 0.725 16.795 1.245 ;
        RECT 12.000 0.110 24.025 0.175 ;
        RECT 21.400 0.110 24.0 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.800 0.535 9.405 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 17.200 0.540 24.09 0.67 ;
        END
    END b
END na02m80

MACRO na02f01
    CLASS CORE ;
    FOREIGN na02f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.450 0.110 0.58 1.215 ;
        RECT 0.430 0.725 0.625 1.245 ;
        RECT 0.450 0.110 0.905 0.175 ;
        RECT 0.805 0.110 0.935 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.070 0.535 0.33 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.645 0.540 0.905 0.67 ;
        END
    END b
END na02f01

MACRO na02f02
    CLASS CORE ;
    FOREIGN na02f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.800 0.110 2.19 1.215 ;
        RECT 1.710 0.725 2.49 1.245 ;
        RECT 1.800 0.110 3.62 0.175 ;
        RECT 3.210 0.110 3.6 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.270 0.535 1.44 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.540 3.62 0.67 ;
        END
    END b
END na02f02

MACRO na02f03
    CLASS CORE ;
    FOREIGN na02f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.250 0.110 2.77 1.215 ;
        RECT 2.140 0.725 3.18 1.245 ;
        RECT 2.250 0.110 4.525 0.175 ;
        RECT 4.015 0.110 4.535 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.340 0.535 1.77 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.225 0.540 4.525 0.67 ;
        END
    END b
END na02f03

MACRO na02f04
    CLASS CORE ;
    FOREIGN na02f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.840 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.700 0.110 3.285 1.215 ;
        RECT 2.565 0.725 3.8 1.245 ;
        RECT 2.700 0.110 5.43 0.175 ;
        RECT 4.815 0.110 5.4 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.405 0.535 2.095 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.870 0.540 5.43 0.67 ;
        END
    END b
END na02f04

MACRO na02f06
    CLASS CORE ;
    FOREIGN na02f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.300 0.110 4.015 1.215 ;
        RECT 3.135 0.725 4.63 1.245 ;
        RECT 3.300 0.110 6.615 0.175 ;
        RECT 5.885 0.110 6.6 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.495 0.535 2.575 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.730 0.540 6.615 0.67 ;
        END
    END b
END na02f06

MACRO na02f08
    CLASS CORE ;
    FOREIGN na02f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.880 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.900 0.110 4.745 1.215 ;
        RECT 3.705 0.725 5.46 1.245 ;
        RECT 3.900 0.110 7.8 0.175 ;
        RECT 6.955 0.110 7.8 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.585 0.535 3.055 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.590 0.540 7.865 0.67 ;
        END
    END b
END na02f08

MACRO na02f10
    CLASS CORE ;
    FOREIGN na02f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.020 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.350 0.110 5.325 1.215 ;
        RECT 4.135 0.725 6.085 1.245 ;
        RECT 4.350 0.110 8.705 0.175 ;
        RECT 7.760 0.110 8.735 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.655 0.535 3.385 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.235 0.540 8.705 0.67 ;
        END
    END b
END na02f10

MACRO na02f20
    CLASS CORE ;
    FOREIGN na02f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.150 0.110 7.515 1.215 ;
        RECT 5.845 0.725 8.64 1.245 ;
        RECT 6.150 0.110 12.325 0.175 ;
        RECT 10.970 0.110 12.335 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.535 4.825 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.815 0.540 12.325 0.67 ;
        END
    END b
END na02f20

MACRO na02f40
    CLASS CORE ;
    FOREIGN na02f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.550 0.110 10.435 1.215 ;
        RECT 8.125 0.725 11.96 1.245 ;
        RECT 8.550 0.110 17.13 0.175 ;
        RECT 15.250 0.110 17.135 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.285 0.535 6.68 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.255 0.540 17.195 0.67 ;
        END
    END b
END na02f40

MACRO na02f80
    CLASS CORE ;
    FOREIGN na02f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.400 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.000 0.110 14.6 1.215 ;
        RECT 11.400 0.725 16.795 1.245 ;
        RECT 12.000 0.110 24.025 0.175 ;
        RECT 21.400 0.110 24.0 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.800 0.535 9.405 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 17.200 0.540 24.09 0.67 ;
        END
    END b
END na02f80

MACRO na03s01
    CLASS CORE ;
    FOREIGN na03s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.555 0.805 0.685 1.26 ;
        RECT 0.555 0.805 1.27 0.87 ;
        RECT 1.165 0.090 1.295 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.050 0.630 0.375 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.470 0.090 0.73 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.850 0.090 1.045 0.74 ;
        END
    END c
END na03s01

MACRO na03s02
    CLASS CORE ;
    FOREIGN na03s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.805 1.65 1.26 ;
        RECT 1.390 0.805 3.145 0.87 ;
        RECT 2.910 0.090 3.17 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.130 0.630 0.91 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.170 0.090 1.885 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.130 0.090 2.65 0.74 ;
        END
    END c
END na03s02

MACRO na03s03
    CLASS CORE ;
    FOREIGN na03s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.805 1.995 1.26 ;
        RECT 1.670 0.805 3.815 0.87 ;
        RECT 3.490 0.090 3.815 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.155 0.630 1.065 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.405 0.090 2.25 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.555 0.090 3.14 0.74 ;
        END
    END c
END na03s03

MACRO na03s04
    CLASS CORE ;
    FOREIGN na03s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.945 0.805 2.335 1.26 ;
        RECT 1.945 0.805 4.415 0.87 ;
        RECT 4.075 0.090 4.465 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.180 0.630 1.22 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.640 0.090 2.615 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.980 0.090 3.695 0.74 ;
        END
    END c
END na03s04

MACRO na03s06
    CLASS CORE ;
    FOREIGN na03s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.365 0.805 2.82 1.26 ;
        RECT 2.365 0.805 5.42 0.87 ;
        RECT 4.945 0.090 5.4 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.220 0.630 1.52 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.990 0.090 3.16 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.620 0.090 4.465 0.74 ;
        END
    END c
END na03s06

MACRO na03s08
    CLASS CORE ;
    FOREIGN na03s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.805 3.3 1.26 ;
        RECT 2.780 0.805 6.355 0.87 ;
        RECT 5.820 0.090 6.34 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.260 0.630 1.755 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.340 0.090 3.77 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.260 0.090 5.235 0.74 ;
        END
    END c
END na03s08

MACRO na03s10
    CLASS CORE ;
    FOREIGN na03s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.060 0.805 3.645 1.26 ;
        RECT 3.060 0.805 6.96 0.87 ;
        RECT 6.400 0.090 6.985 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.285 0.630 1.975 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.575 0.090 4.135 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.685 0.090 5.79 0.74 ;
        END
    END c
END na03s10

MACRO na03s20
    CLASS CORE ;
    FOREIGN na03s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.400 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.170 0.805 4.95 1.26 ;
        RECT 4.170 0.805 9.5 0.87 ;
        RECT 8.730 0.090 9.51 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.390 0.630 2.665 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.510 0.090 5.59 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.390 0.090 7.885 0.74 ;
        END
    END c
END na03s20

MACRO na03s40
    CLASS CORE ;
    FOREIGN na03s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.700 0.805 6.74 1.26 ;
        RECT 5.700 0.805 12.98 0.87 ;
        RECT 11.930 0.090 12.97 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.535 0.630 3.655 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.795 0.090 7.655 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.735 0.090 10.815 0.74 ;
        END
    END c
END na03s40

MACRO na03s80
    CLASS CORE ;
    FOREIGN na03s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.925 0.805 9.42 1.26 ;
        RECT 7.925 0.805 18.065 0.87 ;
        RECT 16.585 0.090 18.08 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.740 0.630 5.095 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.670 0.090 10.635 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.140 0.090 15.0 0.74 ;
        END
    END c
END na03s80

MACRO na03m01
    CLASS CORE ;
    FOREIGN na03m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.555 0.805 0.685 1.26 ;
        RECT 0.555 0.805 1.27 0.87 ;
        RECT 1.165 0.090 1.295 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.050 0.630 0.375 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.470 0.090 0.73 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.850 0.090 1.045 0.74 ;
        END
    END c
END na03m01

MACRO na03m02
    CLASS CORE ;
    FOREIGN na03m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.805 1.65 1.26 ;
        RECT 1.390 0.805 3.145 0.87 ;
        RECT 2.910 0.090 3.17 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.130 0.630 0.91 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.170 0.090 1.885 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.130 0.090 2.65 0.74 ;
        END
    END c
END na03m02

MACRO na03m03
    CLASS CORE ;
    FOREIGN na03m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.805 1.995 1.26 ;
        RECT 1.670 0.805 3.815 0.87 ;
        RECT 3.490 0.090 3.815 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.155 0.630 1.065 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.405 0.090 2.25 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.555 0.090 3.14 0.74 ;
        END
    END c
END na03m03

MACRO na03m04
    CLASS CORE ;
    FOREIGN na03m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.945 0.805 2.335 1.26 ;
        RECT 1.945 0.805 4.415 0.87 ;
        RECT 4.075 0.090 4.465 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.180 0.630 1.22 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.640 0.090 2.615 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.980 0.090 3.695 0.74 ;
        END
    END c
END na03m04

MACRO na03m06
    CLASS CORE ;
    FOREIGN na03m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.365 0.805 2.82 1.26 ;
        RECT 2.365 0.805 5.42 0.87 ;
        RECT 4.945 0.090 5.4 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.220 0.630 1.52 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.990 0.090 3.16 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.620 0.090 4.465 0.74 ;
        END
    END c
END na03m06

MACRO na03m08
    CLASS CORE ;
    FOREIGN na03m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.805 3.3 1.26 ;
        RECT 2.780 0.805 6.355 0.87 ;
        RECT 5.820 0.090 6.34 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.260 0.630 1.755 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.340 0.090 3.77 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.260 0.090 5.235 0.74 ;
        END
    END c
END na03m08

MACRO na03m10
    CLASS CORE ;
    FOREIGN na03m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.060 0.805 3.645 1.26 ;
        RECT 3.060 0.805 6.96 0.87 ;
        RECT 6.400 0.090 6.985 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.285 0.630 1.975 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.575 0.090 4.135 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.685 0.090 5.79 0.74 ;
        END
    END c
END na03m10

MACRO na03m20
    CLASS CORE ;
    FOREIGN na03m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.400 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.170 0.805 4.95 1.26 ;
        RECT 4.170 0.805 9.5 0.87 ;
        RECT 8.730 0.090 9.51 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.390 0.630 2.665 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.510 0.090 5.59 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.390 0.090 7.885 0.74 ;
        END
    END c
END na03m20

MACRO na03m40
    CLASS CORE ;
    FOREIGN na03m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.700 0.805 6.74 1.26 ;
        RECT 5.700 0.805 12.98 0.87 ;
        RECT 11.930 0.090 12.97 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.535 0.630 3.655 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.795 0.090 7.655 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.735 0.090 10.815 0.74 ;
        END
    END c
END na03m40

MACRO na03m80
    CLASS CORE ;
    FOREIGN na03m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.925 0.805 9.42 1.26 ;
        RECT 7.925 0.805 18.065 0.87 ;
        RECT 16.585 0.090 18.08 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.740 0.630 5.095 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.670 0.090 10.635 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.140 0.090 15.0 0.74 ;
        END
    END c
END na03m80

MACRO na03f01
    CLASS CORE ;
    FOREIGN na03f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.555 0.805 0.685 1.26 ;
        RECT 0.555 0.805 1.27 0.87 ;
        RECT 1.165 0.090 1.295 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.050 0.630 0.375 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.470 0.090 0.73 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.850 0.090 1.045 0.74 ;
        END
    END c
END na03f01

MACRO na03f02
    CLASS CORE ;
    FOREIGN na03f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.805 1.65 1.26 ;
        RECT 1.390 0.805 3.145 0.87 ;
        RECT 2.910 0.090 3.17 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.130 0.630 0.91 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.170 0.090 1.885 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.130 0.090 2.65 0.74 ;
        END
    END c
END na03f02

MACRO na03f03
    CLASS CORE ;
    FOREIGN na03f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.805 1.995 1.26 ;
        RECT 1.670 0.805 3.815 0.87 ;
        RECT 3.490 0.090 3.815 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.155 0.630 1.065 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.405 0.090 2.25 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.555 0.090 3.14 0.74 ;
        END
    END c
END na03f03

MACRO na03f04
    CLASS CORE ;
    FOREIGN na03f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.945 0.805 2.335 1.26 ;
        RECT 1.945 0.805 4.415 0.87 ;
        RECT 4.075 0.090 4.465 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.180 0.630 1.22 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.640 0.090 2.615 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.980 0.090 3.695 0.74 ;
        END
    END c
END na03f04

MACRO na03f06
    CLASS CORE ;
    FOREIGN na03f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.365 0.805 2.82 1.26 ;
        RECT 2.365 0.805 5.42 0.87 ;
        RECT 4.945 0.090 5.4 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.220 0.630 1.52 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.990 0.090 3.16 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.620 0.090 4.465 0.74 ;
        END
    END c
END na03f06

MACRO na03f08
    CLASS CORE ;
    FOREIGN na03f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.805 3.3 1.26 ;
        RECT 2.780 0.805 6.355 0.87 ;
        RECT 5.820 0.090 6.34 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.260 0.630 1.755 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.340 0.090 3.77 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.260 0.090 5.235 0.74 ;
        END
    END c
END na03f08

MACRO na03f10
    CLASS CORE ;
    FOREIGN na03f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.060 0.805 3.645 1.26 ;
        RECT 3.060 0.805 6.96 0.87 ;
        RECT 6.400 0.090 6.985 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.285 0.630 1.975 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.575 0.090 4.135 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.685 0.090 5.79 0.74 ;
        END
    END c
END na03f10

MACRO na03f20
    CLASS CORE ;
    FOREIGN na03f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.400 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.170 0.805 4.95 1.26 ;
        RECT 4.170 0.805 9.5 0.87 ;
        RECT 8.730 0.090 9.51 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.390 0.630 2.665 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.510 0.090 5.59 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.390 0.090 7.885 0.74 ;
        END
    END c
END na03f20

MACRO na03f40
    CLASS CORE ;
    FOREIGN na03f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.700 0.805 6.74 1.26 ;
        RECT 5.700 0.805 12.98 0.87 ;
        RECT 11.930 0.090 12.97 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.535 0.630 3.655 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.795 0.090 7.655 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.735 0.090 10.815 0.74 ;
        END
    END c
END na03f40

MACRO na03f80
    CLASS CORE ;
    FOREIGN na03f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.925 0.805 9.42 1.26 ;
        RECT 7.925 0.805 18.065 0.87 ;
        RECT 16.585 0.090 18.08 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.740 0.630 5.095 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.670 0.090 10.635 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.140 0.090 15.0 0.74 ;
        END
    END c
END na03f80

MACRO na04s01
    CLASS CORE ;
    FOREIGN na04s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.210 0.53 0.925 ;
        RECT 0.465 0.870 0.79 0.935 ;
        RECT 0.715 0.870 0.78 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.725 1.34 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.725 1.085 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.635 0.405 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.725 0.83 0.79 ;
        END
    END d
END na04s01

MACRO na04s02
    CLASS CORE ;
    FOREIGN na04s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.180 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.210 1.535 0.925 ;
        RECT 1.275 0.870 2.185 0.935 ;
        RECT 1.970 0.870 2.23 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.145 0.725 3.6 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.445 0.725 2.9 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.580 0.635 1.035 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.750 0.725 2.205 0.79 ;
        END
    END d
END na04s02

MACRO na04s03
    CLASS CORE ;
    FOREIGN na04s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.210 1.945 0.925 ;
        RECT 1.620 0.870 2.79 0.935 ;
        RECT 2.510 0.870 2.835 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.725 4.585 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.725 3.7 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.635 1.32 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.725 2.815 0.79 ;
        END
    END d
END na04s03

MACRO na04s04
    CLASS CORE ;
    FOREIGN na04s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.210 2.18 0.925 ;
        RECT 1.855 0.870 3.22 0.935 ;
        RECT 2.865 0.870 3.19 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.725 5.225 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.725 4.21 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.840 0.635 1.49 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.725 3.195 0.79 ;
        END
    END d
END na04s04

MACRO na04s06
    CLASS CORE ;
    FOREIGN na04s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.220 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.200 0.210 2.59 0.925 ;
        RECT 2.200 0.870 3.825 0.935 ;
        RECT 3.405 0.870 3.795 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.430 0.725 6.21 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.230 0.725 5.01 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.995 0.635 1.775 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.025 0.725 3.805 0.79 ;
        END
    END d
END na04s06

MACRO na04s08
    CLASS CORE ;
    FOREIGN na04s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.550 0.210 3.005 0.925 ;
        RECT 2.550 0.870 4.435 0.935 ;
        RECT 3.940 0.870 4.395 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.290 0.725 7.2 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.895 0.725 5.805 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.155 0.635 2.065 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.500 0.725 4.41 0.79 ;
        END
    END d
END na04s08

MACRO na04s10
    CLASS CORE ;
    FOREIGN na04s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.120 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.210 3.3 0.925 ;
        RECT 2.780 0.870 4.795 0.935 ;
        RECT 4.300 0.870 4.82 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.860 0.725 7.835 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.340 0.725 6.315 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.260 0.635 2.235 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.820 0.725 4.795 0.79 ;
        END
    END d
END na04s10

MACRO na04s20
    CLASS CORE ;
    FOREIGN na04s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.920 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.940 0.210 4.655 0.925 ;
        RECT 3.940 0.870 6.8 0.935 ;
        RECT 6.090 0.870 6.805 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.720 0.725 11.15 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.565 0.725 8.995 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.785 0.635 3.215 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.410 0.725 6.84 0.79 ;
        END
    END d
END na04s20

MACRO na04s40
    CLASS CORE ;
    FOREIGN na04s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.480 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.330 0.210 6.305 0.925 ;
        RECT 5.330 0.870 9.23 0.935 ;
        RECT 8.240 0.870 9.215 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 13.150 0.725 15.035 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.235 0.725 12.12 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.415 0.635 4.3 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.320 0.725 9.205 0.79 ;
        END
    END d
END na04s40

MACRO na04s80
    CLASS CORE ;
    FOREIGN na04s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 24.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.415 0.210 8.78 0.925 ;
        RECT 7.415 0.870 12.875 0.935 ;
        RECT 11.465 0.870 12.83 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 18.295 0.725 20.96 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 14.240 0.725 16.905 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.360 0.635 6.025 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.185 0.725 12.85 0.79 ;
        END
    END d
END na04s80

MACRO na04m01
    CLASS CORE ;
    FOREIGN na04m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.210 0.53 0.925 ;
        RECT 0.465 0.870 0.79 0.935 ;
        RECT 0.715 0.870 0.78 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.725 1.34 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.725 1.085 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.635 0.405 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.725 0.83 0.79 ;
        END
    END d
END na04m01

MACRO na04m02
    CLASS CORE ;
    FOREIGN na04m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.180 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.210 1.535 0.925 ;
        RECT 1.275 0.870 2.185 0.935 ;
        RECT 1.970 0.870 2.23 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.145 0.725 3.6 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.445 0.725 2.9 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.580 0.635 1.035 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.750 0.725 2.205 0.79 ;
        END
    END d
END na04m02

MACRO na04m03
    CLASS CORE ;
    FOREIGN na04m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.210 1.945 0.925 ;
        RECT 1.620 0.870 2.79 0.935 ;
        RECT 2.510 0.870 2.835 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.725 4.585 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.725 3.7 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.635 1.32 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.725 2.815 0.79 ;
        END
    END d
END na04m03

MACRO na04m04
    CLASS CORE ;
    FOREIGN na04m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.210 2.18 0.925 ;
        RECT 1.855 0.870 3.22 0.935 ;
        RECT 2.865 0.870 3.19 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.725 5.225 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.725 4.21 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.840 0.635 1.49 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.725 3.195 0.79 ;
        END
    END d
END na04m04

MACRO na04m06
    CLASS CORE ;
    FOREIGN na04m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.220 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.200 0.210 2.59 0.925 ;
        RECT 2.200 0.870 3.825 0.935 ;
        RECT 3.405 0.870 3.795 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.430 0.725 6.21 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.230 0.725 5.01 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.995 0.635 1.775 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.025 0.725 3.805 0.79 ;
        END
    END d
END na04m06

MACRO na04m08
    CLASS CORE ;
    FOREIGN na04m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.550 0.210 3.005 0.925 ;
        RECT 2.550 0.870 4.435 0.935 ;
        RECT 3.940 0.870 4.395 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.290 0.725 7.2 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.895 0.725 5.805 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.155 0.635 2.065 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.500 0.725 4.41 0.79 ;
        END
    END d
END na04m08

MACRO na04m10
    CLASS CORE ;
    FOREIGN na04m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.120 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.210 3.3 0.925 ;
        RECT 2.780 0.870 4.795 0.935 ;
        RECT 4.300 0.870 4.82 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.860 0.725 7.835 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.340 0.725 6.315 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.260 0.635 2.235 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.820 0.725 4.795 0.79 ;
        END
    END d
END na04m10

MACRO na04m20
    CLASS CORE ;
    FOREIGN na04m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.920 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.940 0.210 4.655 0.925 ;
        RECT 3.940 0.870 6.8 0.935 ;
        RECT 6.090 0.870 6.805 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.720 0.725 11.15 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.565 0.725 8.995 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.785 0.635 3.215 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.410 0.725 6.84 0.79 ;
        END
    END d
END na04m20

MACRO na04m40
    CLASS CORE ;
    FOREIGN na04m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.480 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.330 0.210 6.305 0.925 ;
        RECT 5.330 0.870 9.23 0.935 ;
        RECT 8.240 0.870 9.215 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 13.150 0.725 15.035 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.235 0.725 12.12 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.415 0.635 4.3 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.320 0.725 9.205 0.79 ;
        END
    END d
END na04m40

MACRO na04m80
    CLASS CORE ;
    FOREIGN na04m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 24.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.415 0.210 8.78 0.925 ;
        RECT 7.415 0.870 12.875 0.935 ;
        RECT 11.465 0.870 12.83 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 18.295 0.725 20.96 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 14.240 0.725 16.905 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.360 0.635 6.025 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.185 0.725 12.85 0.79 ;
        END
    END d
END na04m80

MACRO na04f01
    CLASS CORE ;
    FOREIGN na04f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.210 0.53 0.925 ;
        RECT 0.465 0.870 0.79 0.935 ;
        RECT 0.715 0.870 0.78 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.725 1.34 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.725 1.085 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.635 0.405 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.725 0.83 0.79 ;
        END
    END d
END na04f01

MACRO na04f02
    CLASS CORE ;
    FOREIGN na04f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.180 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.210 1.535 0.925 ;
        RECT 1.275 0.870 2.185 0.935 ;
        RECT 1.970 0.870 2.23 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.145 0.725 3.6 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.445 0.725 2.9 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.580 0.635 1.035 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.750 0.725 2.205 0.79 ;
        END
    END d
END na04f02

MACRO na04f03
    CLASS CORE ;
    FOREIGN na04f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.210 1.945 0.925 ;
        RECT 1.620 0.870 2.79 0.935 ;
        RECT 2.510 0.870 2.835 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.725 4.585 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.725 3.7 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.635 1.32 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.725 2.815 0.79 ;
        END
    END d
END na04f03

MACRO na04f04
    CLASS CORE ;
    FOREIGN na04f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.210 2.18 0.925 ;
        RECT 1.855 0.870 3.22 0.935 ;
        RECT 2.865 0.870 3.19 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.725 5.225 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.725 4.21 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.840 0.635 1.49 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.725 3.195 0.79 ;
        END
    END d
END na04f04

MACRO na04f06
    CLASS CORE ;
    FOREIGN na04f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.220 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.200 0.210 2.59 0.925 ;
        RECT 2.200 0.870 3.825 0.935 ;
        RECT 3.405 0.870 3.795 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.430 0.725 6.21 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.230 0.725 5.01 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.995 0.635 1.775 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.025 0.725 3.805 0.79 ;
        END
    END d
END na04f06

MACRO na04f08
    CLASS CORE ;
    FOREIGN na04f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.550 0.210 3.005 0.925 ;
        RECT 2.550 0.870 4.435 0.935 ;
        RECT 3.940 0.870 4.395 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.290 0.725 7.2 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.895 0.725 5.805 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.155 0.635 2.065 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.500 0.725 4.41 0.79 ;
        END
    END d
END na04f08

MACRO na04f10
    CLASS CORE ;
    FOREIGN na04f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.120 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.210 3.3 0.925 ;
        RECT 2.780 0.870 4.795 0.935 ;
        RECT 4.300 0.870 4.82 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.860 0.725 7.835 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.340 0.725 6.315 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.260 0.635 2.235 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.820 0.725 4.795 0.79 ;
        END
    END d
END na04f10

MACRO na04f20
    CLASS CORE ;
    FOREIGN na04f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.920 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.940 0.210 4.655 0.925 ;
        RECT 3.940 0.870 6.8 0.935 ;
        RECT 6.090 0.870 6.805 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.720 0.725 11.15 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.565 0.725 8.995 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.785 0.635 3.215 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.410 0.725 6.84 0.79 ;
        END
    END d
END na04f20

MACRO na04f40
    CLASS CORE ;
    FOREIGN na04f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.480 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.330 0.210 6.305 0.925 ;
        RECT 5.330 0.870 9.23 0.935 ;
        RECT 8.240 0.870 9.215 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 13.150 0.725 15.035 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.235 0.725 12.12 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.415 0.635 4.3 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.320 0.725 9.205 0.79 ;
        END
    END d
END na04f40

MACRO na04f80
    CLASS CORE ;
    FOREIGN na04f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 24.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.415 0.210 8.78 0.925 ;
        RECT 7.415 0.870 12.875 0.935 ;
        RECT 11.465 0.870 12.83 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 18.295 0.725 20.96 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 14.240 0.725 16.905 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.360 0.635 6.025 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.185 0.725 12.85 0.79 ;
        END
    END d
END na04f80

MACRO no02s01
    CLASS CORE ;
    FOREIGN no02s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.520 0.150 0.65 0.54 ;
        RECT 0.465 0.150 0.66 0.28 ;
        RECT 0.520 0.505 0.91 0.57 ;
        RECT 0.805 0.505 0.935 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.235 0.340 0.43 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.715 0.340 0.91 0.405 ;
        END
    END b
END no02s01

MACRO no02s02
    CLASS CORE ;
    FOREIGN no02s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.150 2.475 0.54 ;
        RECT 1.860 0.150 2.64 0.28 ;
        RECT 2.085 0.505 3.58 0.57 ;
        RECT 3.210 0.505 3.6 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.945 0.340 1.725 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.865 0.340 3.645 0.405 ;
        END
    END b
END no02s02

MACRO no02s03
    CLASS CORE ;
    FOREIGN no02s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.605 0.150 3.125 0.54 ;
        RECT 2.325 0.150 3.365 0.28 ;
        RECT 2.605 0.505 4.49 0.57 ;
        RECT 4.015 0.505 4.535 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.180 0.340 2.09 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.580 0.340 4.49 0.405 ;
        END
    END b
END no02s03

MACRO no02s04
    CLASS CORE ;
    FOREIGN no02s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.840 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.130 0.150 3.715 0.54 ;
        RECT 2.790 0.150 4.025 0.28 ;
        RECT 3.130 0.505 5.405 0.57 ;
        RECT 4.815 0.505 5.4 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.420 0.340 2.525 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.340 5.405 0.405 ;
        END
    END b
END no02s04

MACRO no02s06
    CLASS CORE ;
    FOREIGN no02s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.820 0.150 4.535 0.54 ;
        RECT 3.410 0.150 4.905 0.28 ;
        RECT 3.820 0.505 6.615 0.57 ;
        RECT 5.885 0.505 6.6 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.735 0.340 3.1 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.255 0.340 6.62 0.405 ;
        END
    END b
END no02s06

MACRO no02s08
    CLASS CORE ;
    FOREIGN no02s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.880 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.520 0.150 5.365 0.54 ;
        RECT 4.030 0.150 5.785 0.28 ;
        RECT 4.520 0.505 7.835 0.57 ;
        RECT 6.955 0.505 7.8 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.045 0.340 3.67 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.210 0.340 7.835 0.405 ;
        END
    END b
END no02s08

MACRO no02s10
    CLASS CORE ;
    FOREIGN no02s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.020 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.040 0.150 6.015 0.54 ;
        RECT 4.495 0.150 6.445 0.28 ;
        RECT 5.040 0.505 8.68 0.57 ;
        RECT 7.760 0.505 8.735 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.285 0.340 4.105 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.925 0.340 8.745 0.405 ;
        END
    END b
END no02s10

MACRO no02s20
    CLASS CORE ;
    FOREIGN no02s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.125 0.150 8.49 0.54 ;
        RECT 6.355 0.150 9.15 0.28 ;
        RECT 7.125 0.505 12.325 0.57 ;
        RECT 10.970 0.505 12.335 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.230 0.340 5.765 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.790 0.340 12.325 0.405 ;
        END
    END b
END no02s20

MACRO no02s40
    CLASS CORE ;
    FOREIGN no02s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.905 0.150 11.79 0.54 ;
        RECT 8.835 0.150 12.67 0.28 ;
        RECT 9.905 0.505 17.12 0.57 ;
        RECT 15.250 0.505 17.135 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.490 0.340 8.065 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 13.610 0.340 17.185 0.405 ;
        END
    END b
END no02s40

MACRO no02s80
    CLASS CORE ;
    FOREIGN no02s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.400 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 13.900 0.150 16.5 0.54 ;
        RECT 12.400 0.150 17.795 0.28 ;
        RECT 13.900 0.505 23.975 0.57 ;
        RECT 21.400 0.505 24.0 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.300 0.340 11.305 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 19.100 0.340 24.105 0.405 ;
        END
    END b
END no02s80

MACRO no02m01
    CLASS CORE ;
    FOREIGN no02m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.520 0.150 0.65 0.54 ;
        RECT 0.465 0.150 0.66 0.28 ;
        RECT 0.520 0.505 0.91 0.57 ;
        RECT 0.805 0.505 0.935 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.235 0.340 0.43 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.715 0.340 0.91 0.405 ;
        END
    END b
END no02m01

MACRO no02m02
    CLASS CORE ;
    FOREIGN no02m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.150 2.475 0.54 ;
        RECT 1.860 0.150 2.64 0.28 ;
        RECT 2.085 0.505 3.58 0.57 ;
        RECT 3.210 0.505 3.6 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.945 0.340 1.725 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.865 0.340 3.645 0.405 ;
        END
    END b
END no02m02

MACRO no02m03
    CLASS CORE ;
    FOREIGN no02m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.605 0.150 3.125 0.54 ;
        RECT 2.325 0.150 3.365 0.28 ;
        RECT 2.605 0.505 4.49 0.57 ;
        RECT 4.015 0.505 4.535 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.180 0.340 2.09 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.580 0.340 4.49 0.405 ;
        END
    END b
END no02m03

MACRO no02m04
    CLASS CORE ;
    FOREIGN no02m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.840 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.130 0.150 3.715 0.54 ;
        RECT 2.790 0.150 4.025 0.28 ;
        RECT 3.130 0.505 5.405 0.57 ;
        RECT 4.815 0.505 5.4 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.420 0.340 2.525 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.340 5.405 0.405 ;
        END
    END b
END no02m04

MACRO no02m06
    CLASS CORE ;
    FOREIGN no02m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.820 0.150 4.535 0.54 ;
        RECT 3.410 0.150 4.905 0.28 ;
        RECT 3.820 0.505 6.615 0.57 ;
        RECT 5.885 0.505 6.6 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.735 0.340 3.1 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.255 0.340 6.62 0.405 ;
        END
    END b
END no02m06

MACRO no02m08
    CLASS CORE ;
    FOREIGN no02m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.880 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.520 0.150 5.365 0.54 ;
        RECT 4.030 0.150 5.785 0.28 ;
        RECT 4.520 0.505 7.835 0.57 ;
        RECT 6.955 0.505 7.8 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.045 0.340 3.67 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.210 0.340 7.835 0.405 ;
        END
    END b
END no02m08

MACRO no02m10
    CLASS CORE ;
    FOREIGN no02m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.020 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.040 0.150 6.015 0.54 ;
        RECT 4.495 0.150 6.445 0.28 ;
        RECT 5.040 0.505 8.68 0.57 ;
        RECT 7.760 0.505 8.735 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.285 0.340 4.105 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.925 0.340 8.745 0.405 ;
        END
    END b
END no02m10

MACRO no02m20
    CLASS CORE ;
    FOREIGN no02m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.125 0.150 8.49 0.54 ;
        RECT 6.355 0.150 9.15 0.28 ;
        RECT 7.125 0.505 12.325 0.57 ;
        RECT 10.970 0.505 12.335 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.230 0.340 5.765 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.790 0.340 12.325 0.405 ;
        END
    END b
END no02m20

MACRO no02m40
    CLASS CORE ;
    FOREIGN no02m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.905 0.150 11.79 0.54 ;
        RECT 8.835 0.150 12.67 0.28 ;
        RECT 9.905 0.505 17.12 0.57 ;
        RECT 15.250 0.505 17.135 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.490 0.340 8.065 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 13.610 0.340 17.185 0.405 ;
        END
    END b
END no02m40

MACRO no02m80
    CLASS CORE ;
    FOREIGN no02m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.400 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 13.900 0.150 16.5 0.54 ;
        RECT 12.400 0.150 17.795 0.28 ;
        RECT 13.900 0.505 23.975 0.57 ;
        RECT 21.400 0.505 24.0 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.300 0.340 11.305 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 19.100 0.340 24.105 0.405 ;
        END
    END b
END no02m80

MACRO no02f01
    CLASS CORE ;
    FOREIGN no02f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.520 0.150 0.65 0.54 ;
        RECT 0.465 0.150 0.66 0.28 ;
        RECT 0.520 0.505 0.91 0.57 ;
        RECT 0.805 0.505 0.935 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.235 0.340 0.43 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.715 0.340 0.91 0.405 ;
        END
    END b
END no02f01

MACRO no02f02
    CLASS CORE ;
    FOREIGN no02f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.150 2.475 0.54 ;
        RECT 1.860 0.150 2.64 0.28 ;
        RECT 2.085 0.505 3.58 0.57 ;
        RECT 3.210 0.505 3.6 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.945 0.340 1.725 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.865 0.340 3.645 0.405 ;
        END
    END b
END no02f02

MACRO no02f03
    CLASS CORE ;
    FOREIGN no02f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.605 0.150 3.125 0.54 ;
        RECT 2.325 0.150 3.365 0.28 ;
        RECT 2.605 0.505 4.49 0.57 ;
        RECT 4.015 0.505 4.535 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.180 0.340 2.09 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.580 0.340 4.49 0.405 ;
        END
    END b
END no02f03

MACRO no02f04
    CLASS CORE ;
    FOREIGN no02f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.840 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.130 0.150 3.715 0.54 ;
        RECT 2.790 0.150 4.025 0.28 ;
        RECT 3.130 0.505 5.405 0.57 ;
        RECT 4.815 0.505 5.4 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.420 0.340 2.525 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.340 5.405 0.405 ;
        END
    END b
END no02f04

MACRO no02f06
    CLASS CORE ;
    FOREIGN no02f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.820 0.150 4.535 0.54 ;
        RECT 3.410 0.150 4.905 0.28 ;
        RECT 3.820 0.505 6.615 0.57 ;
        RECT 5.885 0.505 6.6 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.735 0.340 3.1 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.255 0.340 6.62 0.405 ;
        END
    END b
END no02f06

MACRO no02f08
    CLASS CORE ;
    FOREIGN no02f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.880 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.520 0.150 5.365 0.54 ;
        RECT 4.030 0.150 5.785 0.28 ;
        RECT 4.520 0.505 7.835 0.57 ;
        RECT 6.955 0.505 7.8 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.045 0.340 3.67 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.210 0.340 7.835 0.405 ;
        END
    END b
END no02f08

MACRO no02f10
    CLASS CORE ;
    FOREIGN no02f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.020 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.040 0.150 6.015 0.54 ;
        RECT 4.495 0.150 6.445 0.28 ;
        RECT 5.040 0.505 8.68 0.57 ;
        RECT 7.760 0.505 8.735 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.285 0.340 4.105 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.925 0.340 8.745 0.405 ;
        END
    END b
END no02f10

MACRO no02f20
    CLASS CORE ;
    FOREIGN no02f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.125 0.150 8.49 0.54 ;
        RECT 6.355 0.150 9.15 0.28 ;
        RECT 7.125 0.505 12.325 0.57 ;
        RECT 10.970 0.505 12.335 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.230 0.340 5.765 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.790 0.340 12.325 0.405 ;
        END
    END b
END no02f20

MACRO no02f40
    CLASS CORE ;
    FOREIGN no02f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.905 0.150 11.79 0.54 ;
        RECT 8.835 0.150 12.67 0.28 ;
        RECT 9.905 0.505 17.12 0.57 ;
        RECT 15.250 0.505 17.135 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.490 0.340 8.065 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 13.610 0.340 17.185 0.405 ;
        END
    END b
END no02f40

MACRO no02f80
    CLASS CORE ;
    FOREIGN no02f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.400 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 13.900 0.150 16.5 0.54 ;
        RECT 12.400 0.150 17.795 0.28 ;
        RECT 13.900 0.505 23.975 0.57 ;
        RECT 21.400 0.505 24.0 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.300 0.340 11.305 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 19.100 0.340 24.105 0.405 ;
        END
    END b
END no02f80

MACRO no03s01
    CLASS CORE ;
    FOREIGN no03s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.560 0.130 0.69 0.39 ;
        RECT 0.560 0.340 1.275 0.405 ;
        RECT 1.160 0.130 1.29 1.625 ;
        RECT 1.160 0.545 1.29 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.110 0.365 0.37 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.555 0.430 0.75 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.860 0.430 1.055 0.56 ;
        END
    END c
END no03s01

MACRO no03s02
    CLASS CORE ;
    FOREIGN no03s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.400 0.130 1.66 0.39 ;
        RECT 1.400 0.340 3.155 0.405 ;
        RECT 2.900 0.130 3.16 1.625 ;
        RECT 2.900 0.545 3.16 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.280 0.365 0.865 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.430 1.845 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.430 2.67 0.56 ;
        END
    END c
END no03s02

MACRO no03s03
    CLASS CORE ;
    FOREIGN no03s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.680 0.130 2.005 0.39 ;
        RECT 1.680 0.340 3.76 0.405 ;
        RECT 3.480 0.130 3.805 1.625 ;
        RECT 3.480 0.545 3.805 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.335 0.365 1.05 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.430 2.255 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.430 3.165 0.56 ;
        END
    END c
END no03s03

MACRO no03s04
    CLASS CORE ;
    FOREIGN no03s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.960 0.130 2.35 0.39 ;
        RECT 1.960 0.340 4.43 0.405 ;
        RECT 4.060 0.130 4.45 1.625 ;
        RECT 4.060 0.545 4.45 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.390 0.365 1.235 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.945 0.430 2.595 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.010 0.430 3.725 0.56 ;
        END
    END c
END no03s04

MACRO no03s06
    CLASS CORE ;
    FOREIGN no03s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.380 0.130 2.835 0.39 ;
        RECT 2.380 0.340 5.37 0.405 ;
        RECT 4.930 0.130 5.385 1.625 ;
        RECT 4.930 0.545 5.385 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.475 0.365 1.515 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.365 0.430 3.145 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.655 0.430 4.5 0.56 ;
        END
    END c
END no03s06

MACRO no03s08
    CLASS CORE ;
    FOREIGN no03s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.800 0.130 3.32 0.39 ;
        RECT 2.800 0.340 6.31 0.405 ;
        RECT 5.800 0.130 6.32 1.625 ;
        RECT 5.800 0.545 6.32 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.560 0.365 1.795 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.430 3.69 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.430 5.275 0.56 ;
        END
    END c
END no03s08

MACRO no03s10
    CLASS CORE ;
    FOREIGN no03s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.080 0.130 3.665 0.39 ;
        RECT 3.080 0.340 6.98 0.405 ;
        RECT 6.380 0.130 6.965 1.625 ;
        RECT 6.380 0.545 6.965 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.615 0.365 1.98 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.060 0.430 4.1 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.730 0.430 5.835 0.56 ;
        END
    END c
END no03s10

MACRO no03s20
    CLASS CORE ;
    FOREIGN no03s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.400 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.200 0.130 4.98 0.39 ;
        RECT 4.200 0.340 9.465 0.405 ;
        RECT 8.700 0.130 9.48 1.625 ;
        RECT 8.700 0.545 9.48 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.840 0.365 2.66 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.170 0.430 5.6 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.450 0.430 7.945 0.56 ;
        END
    END c
END no03s20

MACRO no03s40
    CLASS CORE ;
    FOREIGN no03s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.740 0.130 6.78 0.39 ;
        RECT 5.740 0.340 12.955 0.405 ;
        RECT 11.890 0.130 12.93 1.625 ;
        RECT 11.890 0.545 12.995 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.150 0.365 3.62 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.700 0.430 7.65 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.815 0.430 10.83 0.56 ;
        END
    END c
END no03s40

MACRO no03s80
    CLASS CORE ;
    FOREIGN no03s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.980 0.130 9.475 0.39 ;
        RECT 7.980 0.340 17.99 0.405 ;
        RECT 16.530 0.130 18.025 1.625 ;
        RECT 16.530 0.545 18.09 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.595 0.365 5.04 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.925 0.430 10.59 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.255 0.430 15.05 0.56 ;
        END
    END c
END no03s80

MACRO no03m01
    CLASS CORE ;
    FOREIGN no03m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.560 0.130 0.69 0.39 ;
        RECT 0.560 0.340 1.275 0.405 ;
        RECT 1.160 0.130 1.29 1.625 ;
        RECT 1.160 0.545 1.29 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.110 0.365 0.37 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.555 0.430 0.75 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.860 0.430 1.055 0.56 ;
        END
    END c
END no03m01

MACRO no03m02
    CLASS CORE ;
    FOREIGN no03m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.400 0.130 1.66 0.39 ;
        RECT 1.400 0.340 3.155 0.405 ;
        RECT 2.900 0.130 3.16 1.625 ;
        RECT 2.900 0.545 3.16 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.280 0.365 0.865 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.430 1.845 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.430 2.67 0.56 ;
        END
    END c
END no03m02

MACRO no03m03
    CLASS CORE ;
    FOREIGN no03m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.680 0.130 2.005 0.39 ;
        RECT 1.680 0.340 3.76 0.405 ;
        RECT 3.480 0.130 3.805 1.625 ;
        RECT 3.480 0.545 3.805 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.335 0.365 1.05 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.430 2.255 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.430 3.165 0.56 ;
        END
    END c
END no03m03

MACRO no03m04
    CLASS CORE ;
    FOREIGN no03m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.960 0.130 2.35 0.39 ;
        RECT 1.960 0.340 4.43 0.405 ;
        RECT 4.060 0.130 4.45 1.625 ;
        RECT 4.060 0.545 4.45 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.390 0.365 1.235 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.945 0.430 2.595 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.010 0.430 3.725 0.56 ;
        END
    END c
END no03m04

MACRO no03m06
    CLASS CORE ;
    FOREIGN no03m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.380 0.130 2.835 0.39 ;
        RECT 2.380 0.340 5.37 0.405 ;
        RECT 4.930 0.130 5.385 1.625 ;
        RECT 4.930 0.545 5.385 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.475 0.365 1.515 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.365 0.430 3.145 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.655 0.430 4.5 0.56 ;
        END
    END c
END no03m06

MACRO no03m08
    CLASS CORE ;
    FOREIGN no03m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.800 0.130 3.32 0.39 ;
        RECT 2.800 0.340 6.31 0.405 ;
        RECT 5.800 0.130 6.32 1.625 ;
        RECT 5.800 0.545 6.32 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.560 0.365 1.795 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.430 3.69 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.430 5.275 0.56 ;
        END
    END c
END no03m08

MACRO no03m10
    CLASS CORE ;
    FOREIGN no03m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.080 0.130 3.665 0.39 ;
        RECT 3.080 0.340 6.98 0.405 ;
        RECT 6.380 0.130 6.965 1.625 ;
        RECT 6.380 0.545 6.965 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.615 0.365 1.98 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.060 0.430 4.1 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.730 0.430 5.835 0.56 ;
        END
    END c
END no03m10

MACRO no03m20
    CLASS CORE ;
    FOREIGN no03m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.400 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.200 0.130 4.98 0.39 ;
        RECT 4.200 0.340 9.465 0.405 ;
        RECT 8.700 0.130 9.48 1.625 ;
        RECT 8.700 0.545 9.48 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.840 0.365 2.66 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.170 0.430 5.6 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.450 0.430 7.945 0.56 ;
        END
    END c
END no03m20

MACRO no03m40
    CLASS CORE ;
    FOREIGN no03m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.740 0.130 6.78 0.39 ;
        RECT 5.740 0.340 12.955 0.405 ;
        RECT 11.890 0.130 12.93 1.625 ;
        RECT 11.890 0.545 12.995 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.150 0.365 3.62 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.700 0.430 7.65 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.815 0.430 10.83 0.56 ;
        END
    END c
END no03m40

MACRO no03m80
    CLASS CORE ;
    FOREIGN no03m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.980 0.130 9.475 0.39 ;
        RECT 7.980 0.340 17.99 0.405 ;
        RECT 16.530 0.130 18.025 1.625 ;
        RECT 16.530 0.545 18.09 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.595 0.365 5.04 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.925 0.430 10.59 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.255 0.430 15.05 0.56 ;
        END
    END c
END no03m80

MACRO no03f01
    CLASS CORE ;
    FOREIGN no03f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.560 0.130 0.69 0.39 ;
        RECT 0.560 0.340 1.275 0.405 ;
        RECT 1.160 0.130 1.29 1.625 ;
        RECT 1.160 0.545 1.29 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.110 0.365 0.37 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.555 0.430 0.75 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.860 0.430 1.055 0.56 ;
        END
    END c
END no03f01

MACRO no03f02
    CLASS CORE ;
    FOREIGN no03f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.400 0.130 1.66 0.39 ;
        RECT 1.400 0.340 3.155 0.405 ;
        RECT 2.900 0.130 3.16 1.625 ;
        RECT 2.900 0.545 3.16 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.280 0.365 0.865 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.430 1.845 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.430 2.67 0.56 ;
        END
    END c
END no03f02

MACRO no03f03
    CLASS CORE ;
    FOREIGN no03f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.680 0.130 2.005 0.39 ;
        RECT 1.680 0.340 3.76 0.405 ;
        RECT 3.480 0.130 3.805 1.625 ;
        RECT 3.480 0.545 3.805 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.335 0.365 1.05 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.430 2.255 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.430 3.165 0.56 ;
        END
    END c
END no03f03

MACRO no03f04
    CLASS CORE ;
    FOREIGN no03f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.960 0.130 2.35 0.39 ;
        RECT 1.960 0.340 4.43 0.405 ;
        RECT 4.060 0.130 4.45 1.625 ;
        RECT 4.060 0.545 4.45 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.390 0.365 1.235 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.945 0.430 2.595 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.010 0.430 3.725 0.56 ;
        END
    END c
END no03f04

MACRO no03f06
    CLASS CORE ;
    FOREIGN no03f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.380 0.130 2.835 0.39 ;
        RECT 2.380 0.340 5.37 0.405 ;
        RECT 4.930 0.130 5.385 1.625 ;
        RECT 4.930 0.545 5.385 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.475 0.365 1.515 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.365 0.430 3.145 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.655 0.430 4.5 0.56 ;
        END
    END c
END no03f06

MACRO no03f08
    CLASS CORE ;
    FOREIGN no03f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.800 0.130 3.32 0.39 ;
        RECT 2.800 0.340 6.31 0.405 ;
        RECT 5.800 0.130 6.32 1.625 ;
        RECT 5.800 0.545 6.32 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.560 0.365 1.795 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.430 3.69 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.430 5.275 0.56 ;
        END
    END c
END no03f08

MACRO no03f10
    CLASS CORE ;
    FOREIGN no03f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.080 0.130 3.665 0.39 ;
        RECT 3.080 0.340 6.98 0.405 ;
        RECT 6.380 0.130 6.965 1.625 ;
        RECT 6.380 0.545 6.965 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.615 0.365 1.98 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.060 0.430 4.1 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.730 0.430 5.835 0.56 ;
        END
    END c
END no03f10

MACRO no03f20
    CLASS CORE ;
    FOREIGN no03f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.400 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.200 0.130 4.98 0.39 ;
        RECT 4.200 0.340 9.465 0.405 ;
        RECT 8.700 0.130 9.48 1.625 ;
        RECT 8.700 0.545 9.48 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.840 0.365 2.66 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.170 0.430 5.6 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.450 0.430 7.945 0.56 ;
        END
    END c
END no03f20

MACRO no03f40
    CLASS CORE ;
    FOREIGN no03f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.740 0.130 6.78 0.39 ;
        RECT 5.740 0.340 12.955 0.405 ;
        RECT 11.890 0.130 12.93 1.625 ;
        RECT 11.890 0.545 12.995 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.150 0.365 3.62 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.700 0.430 7.65 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.815 0.430 10.83 0.56 ;
        END
    END c
END no03f40

MACRO no03f80
    CLASS CORE ;
    FOREIGN no03f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.980 0.130 9.475 0.39 ;
        RECT 7.980 0.340 17.99 0.405 ;
        RECT 16.530 0.130 18.025 1.625 ;
        RECT 16.530 0.545 18.09 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.595 0.365 5.04 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.925 0.430 10.59 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.255 0.430 15.05 0.56 ;
        END
    END c
END no03f80

MACRO no04s01
    CLASS CORE ;
    FOREIGN no04s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.090 0.53 1.455 ;
        RECT 0.465 0.090 0.79 0.155 ;
        RECT 0.715 0.090 0.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.530 1.34 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.530 1.085 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.045 0.530 0.305 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.530 0.83 0.66 ;
        END
    END d
END no04s01

MACRO no04s02
    CLASS CORE ;
    FOREIGN no04s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.180 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.090 1.535 1.455 ;
        RECT 1.275 0.090 2.185 0.155 ;
        RECT 1.960 0.090 2.22 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.145 0.530 3.6 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.445 0.530 2.9 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.120 0.530 0.835 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.750 0.530 2.205 0.66 ;
        END
    END d
END no04s02

MACRO no04s03
    CLASS CORE ;
    FOREIGN no04s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.090 1.945 1.455 ;
        RECT 1.620 0.090 2.79 0.155 ;
        RECT 2.495 0.090 2.82 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.530 4.585 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.530 3.7 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.150 0.530 1.06 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.530 2.815 0.66 ;
        END
    END d
END no04s03

MACRO no04s04
    CLASS CORE ;
    FOREIGN no04s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.090 2.18 1.455 ;
        RECT 1.855 0.090 3.22 0.155 ;
        RECT 2.855 0.090 3.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.530 5.225 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.530 4.21 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.175 0.530 1.215 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.530 3.195 0.66 ;
        END
    END d
END no04s04

MACRO no04s06
    CLASS CORE ;
    FOREIGN no04s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.220 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.200 0.090 2.59 1.455 ;
        RECT 2.200 0.090 3.825 0.155 ;
        RECT 3.390 0.090 3.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.430 0.530 6.21 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.230 0.530 5.01 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.205 0.530 1.44 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.025 0.530 3.805 0.66 ;
        END
    END d
END no04s06

MACRO no04s08
    CLASS CORE ;
    FOREIGN no04s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.550 0.090 3.005 1.455 ;
        RECT 2.550 0.090 4.37 0.155 ;
        RECT 3.925 0.090 4.38 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.290 0.530 7.2 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.895 0.530 5.805 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.240 0.530 1.605 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.500 0.530 4.41 0.66 ;
        END
    END d
END no04s08

MACRO no04s10
    CLASS CORE ;
    FOREIGN no04s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.120 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.090 3.3 1.455 ;
        RECT 2.780 0.090 4.795 0.155 ;
        RECT 4.280 0.090 4.8 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.860 0.530 7.835 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.340 0.530 6.315 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.260 0.530 1.755 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.820 0.530 4.795 0.66 ;
        END
    END d
END no04s10

MACRO no04s20
    CLASS CORE ;
    FOREIGN no04s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.920 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.940 0.090 4.655 1.455 ;
        RECT 3.940 0.090 6.8 0.155 ;
        RECT 6.065 0.090 6.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.720 0.530 11.15 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.565 0.530 8.995 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.370 0.530 2.515 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.410 0.530 6.84 0.66 ;
        END
    END d
END no04s20

MACRO no04s40
    CLASS CORE ;
    FOREIGN no04s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.480 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.330 0.090 6.305 1.455 ;
        RECT 5.330 0.090 9.23 0.155 ;
        RECT 8.205 0.090 9.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 13.150 0.530 15.035 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.235 0.530 12.12 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.500 0.530 3.425 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.320 0.530 9.205 0.66 ;
        END
    END d
END no04s40

MACRO no04s80
    CLASS CORE ;
    FOREIGN no04s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 24.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.415 0.090 8.78 1.455 ;
        RECT 7.415 0.090 12.81 0.155 ;
        RECT 11.415 0.090 12.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 18.295 0.530 20.96 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 14.240 0.530 16.905 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.695 0.530 4.725 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.185 0.530 12.85 0.66 ;
        END
    END d
END no04s80

MACRO no04m01
    CLASS CORE ;
    FOREIGN no04m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.090 0.53 1.455 ;
        RECT 0.465 0.090 0.79 0.155 ;
        RECT 0.715 0.090 0.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.530 1.34 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.530 1.085 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.045 0.530 0.305 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.530 0.83 0.66 ;
        END
    END d
END no04m01

MACRO no04m02
    CLASS CORE ;
    FOREIGN no04m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.180 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.090 1.535 1.455 ;
        RECT 1.275 0.090 2.185 0.155 ;
        RECT 1.960 0.090 2.22 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.145 0.530 3.6 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.445 0.530 2.9 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.120 0.530 0.835 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.750 0.530 2.205 0.66 ;
        END
    END d
END no04m02

MACRO no04m03
    CLASS CORE ;
    FOREIGN no04m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.090 1.945 1.455 ;
        RECT 1.620 0.090 2.79 0.155 ;
        RECT 2.495 0.090 2.82 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.530 4.585 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.530 3.7 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.150 0.530 1.06 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.530 2.815 0.66 ;
        END
    END d
END no04m03

MACRO no04m04
    CLASS CORE ;
    FOREIGN no04m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.090 2.18 1.455 ;
        RECT 1.855 0.090 3.22 0.155 ;
        RECT 2.855 0.090 3.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.530 5.225 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.530 4.21 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.175 0.530 1.215 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.530 3.195 0.66 ;
        END
    END d
END no04m04

MACRO no04m06
    CLASS CORE ;
    FOREIGN no04m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.220 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.200 0.090 2.59 1.455 ;
        RECT 2.200 0.090 3.825 0.155 ;
        RECT 3.390 0.090 3.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.430 0.530 6.21 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.230 0.530 5.01 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.205 0.530 1.44 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.025 0.530 3.805 0.66 ;
        END
    END d
END no04m06

MACRO no04m08
    CLASS CORE ;
    FOREIGN no04m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.550 0.090 3.005 1.455 ;
        RECT 2.550 0.090 4.37 0.155 ;
        RECT 3.925 0.090 4.38 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.290 0.530 7.2 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.895 0.530 5.805 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.240 0.530 1.605 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.500 0.530 4.41 0.66 ;
        END
    END d
END no04m08

MACRO no04m10
    CLASS CORE ;
    FOREIGN no04m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.120 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.090 3.3 1.455 ;
        RECT 2.780 0.090 4.795 0.155 ;
        RECT 4.280 0.090 4.8 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.860 0.530 7.835 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.340 0.530 6.315 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.260 0.530 1.755 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.820 0.530 4.795 0.66 ;
        END
    END d
END no04m10

MACRO no04m20
    CLASS CORE ;
    FOREIGN no04m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.920 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.940 0.090 4.655 1.455 ;
        RECT 3.940 0.090 6.8 0.155 ;
        RECT 6.065 0.090 6.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.720 0.530 11.15 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.565 0.530 8.995 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.370 0.530 2.515 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.410 0.530 6.84 0.66 ;
        END
    END d
END no04m20

MACRO no04m40
    CLASS CORE ;
    FOREIGN no04m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.480 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.330 0.090 6.305 1.455 ;
        RECT 5.330 0.090 9.23 0.155 ;
        RECT 8.205 0.090 9.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 13.150 0.530 15.035 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.235 0.530 12.12 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.500 0.530 3.425 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.320 0.530 9.205 0.66 ;
        END
    END d
END no04m40

MACRO no04m80
    CLASS CORE ;
    FOREIGN no04m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 24.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.415 0.090 8.78 1.455 ;
        RECT 7.415 0.090 12.81 0.155 ;
        RECT 11.415 0.090 12.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 18.295 0.530 20.96 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 14.240 0.530 16.905 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.695 0.530 4.725 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.185 0.530 12.85 0.66 ;
        END
    END d
END no04m80

MACRO no04f01
    CLASS CORE ;
    FOREIGN no04f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.090 0.53 1.455 ;
        RECT 0.465 0.090 0.79 0.155 ;
        RECT 0.715 0.090 0.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.530 1.34 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.530 1.085 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.045 0.530 0.305 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.530 0.83 0.66 ;
        END
    END d
END no04f01

MACRO no04f02
    CLASS CORE ;
    FOREIGN no04f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.180 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.090 1.535 1.455 ;
        RECT 1.275 0.090 2.185 0.155 ;
        RECT 1.960 0.090 2.22 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.145 0.530 3.6 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.445 0.530 2.9 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.120 0.530 0.835 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.750 0.530 2.205 0.66 ;
        END
    END d
END no04f02

MACRO no04f03
    CLASS CORE ;
    FOREIGN no04f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.090 1.945 1.455 ;
        RECT 1.620 0.090 2.79 0.155 ;
        RECT 2.495 0.090 2.82 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.530 4.585 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.530 3.7 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.150 0.530 1.06 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.530 2.815 0.66 ;
        END
    END d
END no04f03

MACRO no04f04
    CLASS CORE ;
    FOREIGN no04f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.090 2.18 1.455 ;
        RECT 1.855 0.090 3.22 0.155 ;
        RECT 2.855 0.090 3.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.530 5.225 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.530 4.21 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.175 0.530 1.215 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.530 3.195 0.66 ;
        END
    END d
END no04f04

MACRO no04f06
    CLASS CORE ;
    FOREIGN no04f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.220 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.200 0.090 2.59 1.455 ;
        RECT 2.200 0.090 3.825 0.155 ;
        RECT 3.390 0.090 3.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.430 0.530 6.21 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.230 0.530 5.01 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.205 0.530 1.44 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.025 0.530 3.805 0.66 ;
        END
    END d
END no04f06

MACRO no04f08
    CLASS CORE ;
    FOREIGN no04f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.550 0.090 3.005 1.455 ;
        RECT 2.550 0.090 4.37 0.155 ;
        RECT 3.925 0.090 4.38 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.290 0.530 7.2 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.895 0.530 5.805 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.240 0.530 1.605 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.500 0.530 4.41 0.66 ;
        END
    END d
END no04f08

MACRO no04f10
    CLASS CORE ;
    FOREIGN no04f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.120 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.090 3.3 1.455 ;
        RECT 2.780 0.090 4.795 0.155 ;
        RECT 4.280 0.090 4.8 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.860 0.530 7.835 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.340 0.530 6.315 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.260 0.530 1.755 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.820 0.530 4.795 0.66 ;
        END
    END d
END no04f10

MACRO no04f20
    CLASS CORE ;
    FOREIGN no04f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.920 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.940 0.090 4.655 1.455 ;
        RECT 3.940 0.090 6.8 0.155 ;
        RECT 6.065 0.090 6.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.720 0.530 11.15 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.565 0.530 8.995 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.370 0.530 2.515 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.410 0.530 6.84 0.66 ;
        END
    END d
END no04f20

MACRO no04f40
    CLASS CORE ;
    FOREIGN no04f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.480 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.330 0.090 6.305 1.455 ;
        RECT 5.330 0.090 9.23 0.155 ;
        RECT 8.205 0.090 9.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 13.150 0.530 15.035 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.235 0.530 12.12 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.500 0.530 3.425 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.320 0.530 9.205 0.66 ;
        END
    END d
END no04f40

MACRO no04f80
    CLASS CORE ;
    FOREIGN no04f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 24.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.415 0.090 8.78 1.455 ;
        RECT 7.415 0.090 12.81 0.155 ;
        RECT 11.415 0.090 12.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 18.295 0.530 20.96 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 14.240 0.530 16.905 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.695 0.530 4.725 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.185 0.530 12.85 0.66 ;
        END
    END d
END no04f80

MACRO ao12s01
    CLASS CORE ;
    FOREIGN ao12s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.820 0.100 0.95 0.685 ;
        RECT 0.860 0.635 0.99 0.765 ;
        RECT 0.860 0.750 1.25 0.815 ;
        RECT 1.125 0.750 1.255 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.585 0.445 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.555 0.505 0.685 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.070 0.585 1.265 0.65 ;
        END
    END c
END ao12s01

MACRO ao12s02
    CLASS CORE ;
    FOREIGN ao12s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.050 0.100 2.31 0.685 ;
        RECT 2.150 0.635 2.41 0.765 ;
        RECT 2.150 0.750 3.06 0.815 ;
        RECT 2.810 0.750 3.07 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.585 1.15 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.505 1.78 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.585 3.19 0.65 ;
        END
    END c
END ao12s02

MACRO ao12s03
    CLASS CORE ;
    FOREIGN ao12s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.460 0.100 2.785 0.685 ;
        RECT 2.580 0.635 2.905 0.765 ;
        RECT 2.580 0.750 3.685 0.815 ;
        RECT 3.370 0.750 3.695 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.755 0.585 1.34 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.505 2.125 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.205 0.585 3.79 0.65 ;
        END
    END c
END ao12s03

MACRO ao12s04
    CLASS CORE ;
    FOREIGN ao12s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.870 0.100 3.26 0.685 ;
        RECT 3.010 0.635 3.4 0.765 ;
        RECT 3.010 0.750 4.31 0.815 ;
        RECT 3.935 0.750 4.325 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.880 0.585 1.595 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.945 0.505 2.53 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.740 0.585 4.455 0.65 ;
        END
    END c
END ao12s04

MACRO ao12s06
    CLASS CORE ;
    FOREIGN ao12s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.485 0.100 3.94 0.685 ;
        RECT 3.655 0.635 4.11 0.765 ;
        RECT 3.655 0.750 5.215 0.815 ;
        RECT 4.775 0.750 5.23 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.070 0.585 1.915 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.365 0.505 3.015 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.540 0.585 5.385 0.65 ;
        END
    END c
END ao12s06

MACRO ao12s08
    CLASS CORE ;
    FOREIGN ao12s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.100 0.100 4.62 0.685 ;
        RECT 4.300 0.635 4.82 0.765 ;
        RECT 4.300 0.750 6.12 0.815 ;
        RECT 5.620 0.750 6.14 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.260 0.585 2.235 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.505 3.56 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.340 0.585 6.315 0.65 ;
        END
    END c
END ao12s08

MACRO ao12s10
    CLASS CORE ;
    FOREIGN ao12s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.510 0.100 5.095 0.685 ;
        RECT 4.730 0.635 5.315 0.765 ;
        RECT 4.730 0.750 6.745 0.815 ;
        RECT 6.180 0.750 6.765 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.385 0.585 2.49 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.060 0.505 3.97 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.875 0.585 6.98 0.65 ;
        END
    END c
END ao12s10

MACRO ao12s20
    CLASS CORE ;
    FOREIGN ao12s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.400 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.150 0.100 6.93 0.685 ;
        RECT 6.450 0.635 7.23 0.765 ;
        RECT 6.450 0.750 9.18 0.815 ;
        RECT 8.430 0.750 9.21 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.890 0.585 3.385 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.170 0.505 5.34 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.010 0.585 9.505 0.65 ;
        END
    END c
END ao12s20

MACRO ao12s40
    CLASS CORE ;
    FOREIGN ao12s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.405 0.100 9.445 0.685 ;
        RECT 8.815 0.635 9.855 0.765 ;
        RECT 8.815 0.750 12.585 0.815 ;
        RECT 11.520 0.750 12.56 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.585 0.585 4.665 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.700 0.505 7.325 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.945 0.585 13.025 0.65 ;
        END
    END c
END ao12s40

MACRO ao12s80
    CLASS CORE ;
    FOREIGN ao12s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 11.685 0.100 13.18 0.685 ;
        RECT 12.255 0.635 13.75 0.765 ;
        RECT 12.255 0.750 17.52 0.815 ;
        RECT 16.015 0.750 17.51 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.585 6.45 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.925 0.505 10.2 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 15.220 0.585 18.08 0.65 ;
        END
    END c
END ao12s80

MACRO ao12m01
    CLASS CORE ;
    FOREIGN ao12m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.820 0.100 0.95 0.685 ;
        RECT 0.860 0.635 0.99 0.765 ;
        RECT 0.860 0.750 1.25 0.815 ;
        RECT 1.125 0.750 1.255 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.585 0.445 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.555 0.505 0.685 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.070 0.585 1.265 0.65 ;
        END
    END c
END ao12m01

MACRO ao12m02
    CLASS CORE ;
    FOREIGN ao12m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.050 0.100 2.31 0.685 ;
        RECT 2.150 0.635 2.41 0.765 ;
        RECT 2.150 0.750 3.06 0.815 ;
        RECT 2.810 0.750 3.07 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.585 1.15 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.505 1.78 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.585 3.19 0.65 ;
        END
    END c
END ao12m02

MACRO ao12m03
    CLASS CORE ;
    FOREIGN ao12m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.460 0.100 2.785 0.685 ;
        RECT 2.580 0.635 2.905 0.765 ;
        RECT 2.580 0.750 3.685 0.815 ;
        RECT 3.370 0.750 3.695 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.755 0.585 1.34 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.505 2.125 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.205 0.585 3.79 0.65 ;
        END
    END c
END ao12m03

MACRO ao12m04
    CLASS CORE ;
    FOREIGN ao12m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.870 0.100 3.26 0.685 ;
        RECT 3.010 0.635 3.4 0.765 ;
        RECT 3.010 0.750 4.31 0.815 ;
        RECT 3.935 0.750 4.325 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.880 0.585 1.595 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.945 0.505 2.53 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.740 0.585 4.455 0.65 ;
        END
    END c
END ao12m04

MACRO ao12m06
    CLASS CORE ;
    FOREIGN ao12m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.485 0.100 3.94 0.685 ;
        RECT 3.655 0.635 4.11 0.765 ;
        RECT 3.655 0.750 5.215 0.815 ;
        RECT 4.775 0.750 5.23 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.070 0.585 1.915 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.365 0.505 3.015 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.540 0.585 5.385 0.65 ;
        END
    END c
END ao12m06

MACRO ao12m08
    CLASS CORE ;
    FOREIGN ao12m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.100 0.100 4.62 0.685 ;
        RECT 4.300 0.635 4.82 0.765 ;
        RECT 4.300 0.750 6.12 0.815 ;
        RECT 5.620 0.750 6.14 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.260 0.585 2.235 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.505 3.56 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.340 0.585 6.315 0.65 ;
        END
    END c
END ao12m08

MACRO ao12m10
    CLASS CORE ;
    FOREIGN ao12m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.510 0.100 5.095 0.685 ;
        RECT 4.730 0.635 5.315 0.765 ;
        RECT 4.730 0.750 6.745 0.815 ;
        RECT 6.180 0.750 6.765 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.385 0.585 2.49 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.060 0.505 3.97 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.875 0.585 6.98 0.65 ;
        END
    END c
END ao12m10

MACRO ao12m20
    CLASS CORE ;
    FOREIGN ao12m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.400 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.150 0.100 6.93 0.685 ;
        RECT 6.450 0.635 7.23 0.765 ;
        RECT 6.450 0.750 9.18 0.815 ;
        RECT 8.430 0.750 9.21 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.890 0.585 3.385 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.170 0.505 5.34 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.010 0.585 9.505 0.65 ;
        END
    END c
END ao12m20

MACRO ao12m40
    CLASS CORE ;
    FOREIGN ao12m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.405 0.100 9.445 0.685 ;
        RECT 8.815 0.635 9.855 0.765 ;
        RECT 8.815 0.750 12.585 0.815 ;
        RECT 11.520 0.750 12.56 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.585 0.585 4.665 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.700 0.505 7.325 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.945 0.585 13.025 0.65 ;
        END
    END c
END ao12m40

MACRO ao12m80
    CLASS CORE ;
    FOREIGN ao12m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 11.685 0.100 13.18 0.685 ;
        RECT 12.255 0.635 13.75 0.765 ;
        RECT 12.255 0.750 17.52 0.815 ;
        RECT 16.015 0.750 17.51 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.585 6.45 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.925 0.505 10.2 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 15.220 0.585 18.08 0.65 ;
        END
    END c
END ao12m80

MACRO ao12f01
    CLASS CORE ;
    FOREIGN ao12f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.820 0.100 0.95 0.685 ;
        RECT 0.860 0.635 0.99 0.765 ;
        RECT 0.860 0.750 1.25 0.815 ;
        RECT 1.125 0.750 1.255 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.585 0.445 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.555 0.505 0.685 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.070 0.585 1.265 0.65 ;
        END
    END c
END ao12f01

MACRO ao12f02
    CLASS CORE ;
    FOREIGN ao12f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.050 0.100 2.31 0.685 ;
        RECT 2.150 0.635 2.41 0.765 ;
        RECT 2.150 0.750 3.06 0.815 ;
        RECT 2.810 0.750 3.07 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.585 1.15 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.505 1.78 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.585 3.19 0.65 ;
        END
    END c
END ao12f02

MACRO ao12f03
    CLASS CORE ;
    FOREIGN ao12f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.460 0.100 2.785 0.685 ;
        RECT 2.580 0.635 2.905 0.765 ;
        RECT 2.580 0.750 3.685 0.815 ;
        RECT 3.370 0.750 3.695 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.755 0.585 1.34 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.505 2.125 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.205 0.585 3.79 0.65 ;
        END
    END c
END ao12f03

MACRO ao12f04
    CLASS CORE ;
    FOREIGN ao12f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.870 0.100 3.26 0.685 ;
        RECT 3.010 0.635 3.4 0.765 ;
        RECT 3.010 0.750 4.31 0.815 ;
        RECT 3.935 0.750 4.325 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.880 0.585 1.595 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.945 0.505 2.53 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.740 0.585 4.455 0.65 ;
        END
    END c
END ao12f04

MACRO ao12f06
    CLASS CORE ;
    FOREIGN ao12f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.485 0.100 3.94 0.685 ;
        RECT 3.655 0.635 4.11 0.765 ;
        RECT 3.655 0.750 5.215 0.815 ;
        RECT 4.775 0.750 5.23 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.070 0.585 1.915 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.365 0.505 3.015 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.540 0.585 5.385 0.65 ;
        END
    END c
END ao12f06

MACRO ao12f08
    CLASS CORE ;
    FOREIGN ao12f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.100 0.100 4.62 0.685 ;
        RECT 4.300 0.635 4.82 0.765 ;
        RECT 4.300 0.750 6.12 0.815 ;
        RECT 5.620 0.750 6.14 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.260 0.585 2.235 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.505 3.56 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.340 0.585 6.315 0.65 ;
        END
    END c
END ao12f08

MACRO ao12f10
    CLASS CORE ;
    FOREIGN ao12f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.510 0.100 5.095 0.685 ;
        RECT 4.730 0.635 5.315 0.765 ;
        RECT 4.730 0.750 6.745 0.815 ;
        RECT 6.180 0.750 6.765 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.385 0.585 2.49 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.060 0.505 3.97 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.875 0.585 6.98 0.65 ;
        END
    END c
END ao12f10

MACRO ao12f20
    CLASS CORE ;
    FOREIGN ao12f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.400 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.150 0.100 6.93 0.685 ;
        RECT 6.450 0.635 7.23 0.765 ;
        RECT 6.450 0.750 9.18 0.815 ;
        RECT 8.430 0.750 9.21 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.890 0.585 3.385 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.170 0.505 5.34 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.010 0.585 9.505 0.65 ;
        END
    END c
END ao12f20

MACRO ao12f40
    CLASS CORE ;
    FOREIGN ao12f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.405 0.100 9.445 0.685 ;
        RECT 8.815 0.635 9.855 0.765 ;
        RECT 8.815 0.750 12.585 0.815 ;
        RECT 11.520 0.750 12.56 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.585 0.585 4.665 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.700 0.505 7.325 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.945 0.585 13.025 0.65 ;
        END
    END c
END ao12f40

MACRO ao12f80
    CLASS CORE ;
    FOREIGN ao12f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 11.685 0.100 13.18 0.685 ;
        RECT 12.255 0.635 13.75 0.765 ;
        RECT 12.255 0.750 17.52 0.815 ;
        RECT 16.015 0.750 17.51 1.53 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.585 6.45 0.65 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.925 0.505 10.2 0.57 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 15.220 0.585 18.08 0.65 ;
        END
    END c
END ao12f80

MACRO ao22s01
    CLASS CORE ;
    FOREIGN ao22s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.090 0.53 1.455 ;
        RECT 0.465 0.090 0.79 0.155 ;
        RECT 0.715 0.090 0.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.530 1.34 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.530 1.085 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.045 0.530 0.305 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.530 0.83 0.66 ;
        END
    END d
END ao22s01

MACRO ao22s02
    CLASS CORE ;
    FOREIGN ao22s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.180 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.090 1.535 1.455 ;
        RECT 1.275 0.090 2.185 0.155 ;
        RECT 1.960 0.090 2.22 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.145 0.530 3.6 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.445 0.530 2.9 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.120 0.530 0.835 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.750 0.530 2.205 0.66 ;
        END
    END d
END ao22s02

MACRO ao22s03
    CLASS CORE ;
    FOREIGN ao22s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.090 1.945 1.455 ;
        RECT 1.620 0.090 2.79 0.155 ;
        RECT 2.495 0.090 2.82 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.530 4.585 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.530 3.7 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.150 0.530 1.06 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.530 2.815 0.66 ;
        END
    END d
END ao22s03

MACRO ao22s04
    CLASS CORE ;
    FOREIGN ao22s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.090 2.18 1.455 ;
        RECT 1.855 0.090 3.22 0.155 ;
        RECT 2.855 0.090 3.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.530 5.225 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.530 4.21 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.175 0.530 1.215 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.530 3.195 0.66 ;
        END
    END d
END ao22s04

MACRO ao22s06
    CLASS CORE ;
    FOREIGN ao22s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.220 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.200 0.090 2.59 1.455 ;
        RECT 2.200 0.090 3.825 0.155 ;
        RECT 3.390 0.090 3.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.430 0.530 6.21 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.230 0.530 5.01 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.205 0.530 1.44 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.025 0.530 3.805 0.66 ;
        END
    END d
END ao22s06

MACRO ao22s08
    CLASS CORE ;
    FOREIGN ao22s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.550 0.090 3.005 1.455 ;
        RECT 2.550 0.090 4.37 0.155 ;
        RECT 3.925 0.090 4.38 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.290 0.530 7.2 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.895 0.530 5.805 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.240 0.530 1.605 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.500 0.530 4.41 0.66 ;
        END
    END d
END ao22s08

MACRO ao22s10
    CLASS CORE ;
    FOREIGN ao22s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.120 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.090 3.3 1.455 ;
        RECT 2.780 0.090 4.795 0.155 ;
        RECT 4.280 0.090 4.8 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.860 0.530 7.835 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.340 0.530 6.315 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.260 0.530 1.755 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.820 0.530 4.795 0.66 ;
        END
    END d
END ao22s10

MACRO ao22s20
    CLASS CORE ;
    FOREIGN ao22s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.920 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.940 0.090 4.655 1.455 ;
        RECT 3.940 0.090 6.8 0.155 ;
        RECT 6.065 0.090 6.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.720 0.530 11.15 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.565 0.530 8.995 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.370 0.530 2.515 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.410 0.530 6.84 0.66 ;
        END
    END d
END ao22s20

MACRO ao22s40
    CLASS CORE ;
    FOREIGN ao22s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.480 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.330 0.090 6.305 1.455 ;
        RECT 5.330 0.090 9.23 0.155 ;
        RECT 8.205 0.090 9.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 13.150 0.530 15.035 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.235 0.530 12.12 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.500 0.530 3.425 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.320 0.530 9.205 0.66 ;
        END
    END d
END ao22s40

MACRO ao22s80
    CLASS CORE ;
    FOREIGN ao22s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 24.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.415 0.090 8.78 1.455 ;
        RECT 7.415 0.090 12.81 0.155 ;
        RECT 11.415 0.090 12.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 18.295 0.530 20.96 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 14.240 0.530 16.905 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.695 0.530 4.725 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.185 0.530 12.85 0.66 ;
        END
    END d
END ao22s80

MACRO ao22m01
    CLASS CORE ;
    FOREIGN ao22m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.090 0.53 1.455 ;
        RECT 0.465 0.090 0.79 0.155 ;
        RECT 0.715 0.090 0.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.530 1.34 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.530 1.085 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.045 0.530 0.305 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.530 0.83 0.66 ;
        END
    END d
END ao22m01

MACRO ao22m02
    CLASS CORE ;
    FOREIGN ao22m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.180 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.090 1.535 1.455 ;
        RECT 1.275 0.090 2.185 0.155 ;
        RECT 1.960 0.090 2.22 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.145 0.530 3.6 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.445 0.530 2.9 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.120 0.530 0.835 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.750 0.530 2.205 0.66 ;
        END
    END d
END ao22m02

MACRO ao22m03
    CLASS CORE ;
    FOREIGN ao22m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.090 1.945 1.455 ;
        RECT 1.620 0.090 2.79 0.155 ;
        RECT 2.495 0.090 2.82 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.530 4.585 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.530 3.7 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.150 0.530 1.06 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.530 2.815 0.66 ;
        END
    END d
END ao22m03

MACRO ao22m04
    CLASS CORE ;
    FOREIGN ao22m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.090 2.18 1.455 ;
        RECT 1.855 0.090 3.22 0.155 ;
        RECT 2.855 0.090 3.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.530 5.225 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.530 4.21 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.175 0.530 1.215 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.530 3.195 0.66 ;
        END
    END d
END ao22m04

MACRO ao22m06
    CLASS CORE ;
    FOREIGN ao22m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.220 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.200 0.090 2.59 1.455 ;
        RECT 2.200 0.090 3.825 0.155 ;
        RECT 3.390 0.090 3.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.430 0.530 6.21 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.230 0.530 5.01 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.205 0.530 1.44 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.025 0.530 3.805 0.66 ;
        END
    END d
END ao22m06

MACRO ao22m08
    CLASS CORE ;
    FOREIGN ao22m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.550 0.090 3.005 1.455 ;
        RECT 2.550 0.090 4.37 0.155 ;
        RECT 3.925 0.090 4.38 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.290 0.530 7.2 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.895 0.530 5.805 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.240 0.530 1.605 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.500 0.530 4.41 0.66 ;
        END
    END d
END ao22m08

MACRO ao22m10
    CLASS CORE ;
    FOREIGN ao22m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.120 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.090 3.3 1.455 ;
        RECT 2.780 0.090 4.795 0.155 ;
        RECT 4.280 0.090 4.8 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.860 0.530 7.835 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.340 0.530 6.315 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.260 0.530 1.755 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.820 0.530 4.795 0.66 ;
        END
    END d
END ao22m10

MACRO ao22m20
    CLASS CORE ;
    FOREIGN ao22m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.920 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.940 0.090 4.655 1.455 ;
        RECT 3.940 0.090 6.8 0.155 ;
        RECT 6.065 0.090 6.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.720 0.530 11.15 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.565 0.530 8.995 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.370 0.530 2.515 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.410 0.530 6.84 0.66 ;
        END
    END d
END ao22m20

MACRO ao22m40
    CLASS CORE ;
    FOREIGN ao22m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.480 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.330 0.090 6.305 1.455 ;
        RECT 5.330 0.090 9.23 0.155 ;
        RECT 8.205 0.090 9.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 13.150 0.530 15.035 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.235 0.530 12.12 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.500 0.530 3.425 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.320 0.530 9.205 0.66 ;
        END
    END d
END ao22m40

MACRO ao22m80
    CLASS CORE ;
    FOREIGN ao22m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 24.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.415 0.090 8.78 1.455 ;
        RECT 7.415 0.090 12.81 0.155 ;
        RECT 11.415 0.090 12.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 18.295 0.530 20.96 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 14.240 0.530 16.905 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.695 0.530 4.725 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.185 0.530 12.85 0.66 ;
        END
    END d
END ao22m80

MACRO ao22f01
    CLASS CORE ;
    FOREIGN ao22f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.090 0.53 1.455 ;
        RECT 0.465 0.090 0.79 0.155 ;
        RECT 0.715 0.090 0.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.530 1.34 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.530 1.085 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.045 0.530 0.305 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.530 0.83 0.66 ;
        END
    END d
END ao22f01

MACRO ao22f02
    CLASS CORE ;
    FOREIGN ao22f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.180 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.090 1.535 1.455 ;
        RECT 1.275 0.090 2.185 0.155 ;
        RECT 1.960 0.090 2.22 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.145 0.530 3.6 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.445 0.530 2.9 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.120 0.530 0.835 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.750 0.530 2.205 0.66 ;
        END
    END d
END ao22f02

MACRO ao22f03
    CLASS CORE ;
    FOREIGN ao22f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.090 1.945 1.455 ;
        RECT 1.620 0.090 2.79 0.155 ;
        RECT 2.495 0.090 2.82 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.530 4.585 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.530 3.7 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.150 0.530 1.06 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.530 2.815 0.66 ;
        END
    END d
END ao22f03

MACRO ao22f04
    CLASS CORE ;
    FOREIGN ao22f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.090 2.18 1.455 ;
        RECT 1.855 0.090 3.22 0.155 ;
        RECT 2.855 0.090 3.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.530 5.225 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.530 4.21 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.175 0.530 1.215 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.530 3.195 0.66 ;
        END
    END d
END ao22f04

MACRO ao22f06
    CLASS CORE ;
    FOREIGN ao22f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.220 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.200 0.090 2.59 1.455 ;
        RECT 2.200 0.090 3.825 0.155 ;
        RECT 3.390 0.090 3.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.430 0.530 6.21 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.230 0.530 5.01 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.205 0.530 1.44 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.025 0.530 3.805 0.66 ;
        END
    END d
END ao22f06

MACRO ao22f08
    CLASS CORE ;
    FOREIGN ao22f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.550 0.090 3.005 1.455 ;
        RECT 2.550 0.090 4.37 0.155 ;
        RECT 3.925 0.090 4.38 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.290 0.530 7.2 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.895 0.530 5.805 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.240 0.530 1.605 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.500 0.530 4.41 0.66 ;
        END
    END d
END ao22f08

MACRO ao22f10
    CLASS CORE ;
    FOREIGN ao22f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.120 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.090 3.3 1.455 ;
        RECT 2.780 0.090 4.795 0.155 ;
        RECT 4.280 0.090 4.8 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.860 0.530 7.835 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.340 0.530 6.315 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.260 0.530 1.755 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.820 0.530 4.795 0.66 ;
        END
    END d
END ao22f10

MACRO ao22f20
    CLASS CORE ;
    FOREIGN ao22f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.920 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.940 0.090 4.655 1.455 ;
        RECT 3.940 0.090 6.8 0.155 ;
        RECT 6.065 0.090 6.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.720 0.530 11.15 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.565 0.530 8.995 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.370 0.530 2.515 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.410 0.530 6.84 0.66 ;
        END
    END d
END ao22f20

MACRO ao22f40
    CLASS CORE ;
    FOREIGN ao22f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.480 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.330 0.090 6.305 1.455 ;
        RECT 5.330 0.090 9.23 0.155 ;
        RECT 8.205 0.090 9.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 13.150 0.530 15.035 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.235 0.530 12.12 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.500 0.530 3.425 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.320 0.530 9.205 0.66 ;
        END
    END d
END ao22f40

MACRO ao22f80
    CLASS CORE ;
    FOREIGN ao22f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 24.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.415 0.090 8.78 1.455 ;
        RECT 7.415 0.090 12.81 0.155 ;
        RECT 11.415 0.090 12.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 18.295 0.530 20.96 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 14.240 0.530 16.905 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.695 0.530 4.725 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.185 0.530 12.85 0.66 ;
        END
    END d
END ao22f80

MACRO oa12s01
    CLASS CORE ;
    FOREIGN oa12s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.860 0.650 0.99 1.235 ;
        RECT 0.750 0.900 0.945 1.225 ;
        RECT 1.100 0.135 1.23 0.72 ;
        RECT 0.860 0.650 1.185 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.720 0.445 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.555 0.720 0.685 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.070 0.740 1.265 0.805 ;
        END
    END c
END oa12s01

MACRO oa12s02
    CLASS CORE ;
    FOREIGN oa12s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.650 2.41 1.235 ;
        RECT 1.870 0.900 2.39 1.225 ;
        RECT 2.750 0.135 3.01 0.72 ;
        RECT 2.150 0.650 2.995 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.720 1.085 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.720 1.715 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.740 3.19 0.805 ;
        END
    END c
END oa12s02

MACRO oa12s03
    CLASS CORE ;
    FOREIGN oa12s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.650 2.905 1.235 ;
        RECT 2.245 0.900 2.895 1.225 ;
        RECT 3.300 0.135 3.625 0.72 ;
        RECT 2.580 0.650 3.62 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.755 0.720 1.275 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.720 2.06 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.205 0.740 3.79 0.805 ;
        END
    END c
END oa12s03

MACRO oa12s04
    CLASS CORE ;
    FOREIGN oa12s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.010 0.650 3.4 1.235 ;
        RECT 2.620 0.900 3.4 1.225 ;
        RECT 3.850 0.135 4.24 0.72 ;
        RECT 3.010 0.650 4.245 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.880 0.720 1.465 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.945 0.720 2.4 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.740 0.740 4.455 0.805 ;
        END
    END c
END oa12s04

MACRO oa12s06
    CLASS CORE ;
    FOREIGN oa12s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.655 0.650 4.11 1.235 ;
        RECT 3.180 0.900 4.09 1.225 ;
        RECT 4.675 0.135 5.13 0.72 ;
        RECT 3.655 0.650 5.085 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.070 0.720 1.85 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.365 0.720 2.885 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.540 0.740 5.385 0.805 ;
        END
    END c
END oa12s06

MACRO oa12s08
    CLASS CORE ;
    FOREIGN oa12s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.650 4.82 1.235 ;
        RECT 3.740 0.900 4.845 1.225 ;
        RECT 5.500 0.135 6.02 0.72 ;
        RECT 4.300 0.650 5.99 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.260 0.720 2.17 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.720 3.43 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.340 0.740 6.315 0.805 ;
        END
    END c
END oa12s08

MACRO oa12s10
    CLASS CORE ;
    FOREIGN oa12s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.730 0.650 5.315 1.235 ;
        RECT 4.115 0.900 5.285 1.225 ;
        RECT 6.050 0.135 6.635 0.72 ;
        RECT 4.730 0.650 6.615 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.385 0.720 2.36 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.060 0.720 3.775 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.875 0.740 6.98 0.805 ;
        END
    END c
END oa12s10

MACRO oa12s20
    CLASS CORE ;
    FOREIGN oa12s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.400 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.450 0.650 7.23 1.235 ;
        RECT 5.610 0.900 7.235 1.225 ;
        RECT 8.250 0.135 9.03 0.72 ;
        RECT 6.450 0.650 9.05 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.890 0.720 3.19 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.170 0.720 5.145 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.010 0.740 9.505 0.805 ;
        END
    END c
END oa12s20

MACRO oa12s40
    CLASS CORE ;
    FOREIGN oa12s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.815 0.650 9.855 1.235 ;
        RECT 7.665 0.900 9.875 1.225 ;
        RECT 11.275 0.135 12.315 0.72 ;
        RECT 8.815 0.650 12.325 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.585 0.720 4.405 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.700 0.720 7.0 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.945 0.740 13.025 0.805 ;
        END
    END c
END oa12s40

MACRO oa12s80
    CLASS CORE ;
    FOREIGN oa12s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.255 0.650 13.75 1.235 ;
        RECT 10.660 0.900 13.715 1.225 ;
        RECT 15.675 0.135 17.17 0.72 ;
        RECT 12.255 0.650 17.13 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.720 6.125 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.925 0.720 9.745 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 15.220 0.740 18.08 0.805 ;
        END
    END c
END oa12s80

MACRO oa12m01
    CLASS CORE ;
    FOREIGN oa12m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.860 0.650 0.99 1.235 ;
        RECT 0.750 0.900 0.945 1.225 ;
        RECT 1.100 0.135 1.23 0.72 ;
        RECT 0.860 0.650 1.185 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.720 0.445 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.555 0.720 0.685 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.070 0.740 1.265 0.805 ;
        END
    END c
END oa12m01

MACRO oa12m02
    CLASS CORE ;
    FOREIGN oa12m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.650 2.41 1.235 ;
        RECT 1.870 0.900 2.39 1.225 ;
        RECT 2.750 0.135 3.01 0.72 ;
        RECT 2.150 0.650 2.995 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.720 1.085 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.720 1.715 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.740 3.19 0.805 ;
        END
    END c
END oa12m02

MACRO oa12m03
    CLASS CORE ;
    FOREIGN oa12m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.650 2.905 1.235 ;
        RECT 2.245 0.900 2.895 1.225 ;
        RECT 3.300 0.135 3.625 0.72 ;
        RECT 2.580 0.650 3.62 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.755 0.720 1.275 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.720 2.06 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.205 0.740 3.79 0.805 ;
        END
    END c
END oa12m03

MACRO oa12m04
    CLASS CORE ;
    FOREIGN oa12m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.010 0.650 3.4 1.235 ;
        RECT 2.620 0.900 3.4 1.225 ;
        RECT 3.850 0.135 4.24 0.72 ;
        RECT 3.010 0.650 4.245 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.880 0.720 1.465 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.945 0.720 2.4 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.740 0.740 4.455 0.805 ;
        END
    END c
END oa12m04

MACRO oa12m06
    CLASS CORE ;
    FOREIGN oa12m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.655 0.650 4.11 1.235 ;
        RECT 3.180 0.900 4.09 1.225 ;
        RECT 4.675 0.135 5.13 0.72 ;
        RECT 3.655 0.650 5.085 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.070 0.720 1.85 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.365 0.720 2.885 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.540 0.740 5.385 0.805 ;
        END
    END c
END oa12m06

MACRO oa12m08
    CLASS CORE ;
    FOREIGN oa12m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.650 4.82 1.235 ;
        RECT 3.740 0.900 4.845 1.225 ;
        RECT 5.500 0.135 6.02 0.72 ;
        RECT 4.300 0.650 5.99 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.260 0.720 2.17 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.720 3.43 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.340 0.740 6.315 0.805 ;
        END
    END c
END oa12m08

MACRO oa12m10
    CLASS CORE ;
    FOREIGN oa12m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.730 0.650 5.315 1.235 ;
        RECT 4.115 0.900 5.285 1.225 ;
        RECT 6.050 0.135 6.635 0.72 ;
        RECT 4.730 0.650 6.615 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.385 0.720 2.36 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.060 0.720 3.775 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.875 0.740 6.98 0.805 ;
        END
    END c
END oa12m10

MACRO oa12m20
    CLASS CORE ;
    FOREIGN oa12m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.400 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.450 0.650 7.23 1.235 ;
        RECT 5.610 0.900 7.235 1.225 ;
        RECT 8.250 0.135 9.03 0.72 ;
        RECT 6.450 0.650 9.05 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.890 0.720 3.19 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.170 0.720 5.145 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.010 0.740 9.505 0.805 ;
        END
    END c
END oa12m20

MACRO oa12m40
    CLASS CORE ;
    FOREIGN oa12m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.815 0.650 9.855 1.235 ;
        RECT 7.665 0.900 9.875 1.225 ;
        RECT 11.275 0.135 12.315 0.72 ;
        RECT 8.815 0.650 12.325 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.585 0.720 4.405 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.700 0.720 7.0 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.945 0.740 13.025 0.805 ;
        END
    END c
END oa12m40

MACRO oa12m80
    CLASS CORE ;
    FOREIGN oa12m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.255 0.650 13.75 1.235 ;
        RECT 10.660 0.900 13.715 1.225 ;
        RECT 15.675 0.135 17.17 0.72 ;
        RECT 12.255 0.650 17.13 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.720 6.125 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.925 0.720 9.745 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 15.220 0.740 18.08 0.805 ;
        END
    END c
END oa12m80

MACRO oa12f01
    CLASS CORE ;
    FOREIGN oa12f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.860 0.650 0.99 1.235 ;
        RECT 0.750 0.900 0.945 1.225 ;
        RECT 1.100 0.135 1.23 0.72 ;
        RECT 0.860 0.650 1.185 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.720 0.445 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.555 0.720 0.685 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.070 0.740 1.265 0.805 ;
        END
    END c
END oa12f01

MACRO oa12f02
    CLASS CORE ;
    FOREIGN oa12f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.650 2.41 1.235 ;
        RECT 1.870 0.900 2.39 1.225 ;
        RECT 2.750 0.135 3.01 0.72 ;
        RECT 2.150 0.650 2.995 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.720 1.085 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.720 1.715 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.740 3.19 0.805 ;
        END
    END c
END oa12f02

MACRO oa12f03
    CLASS CORE ;
    FOREIGN oa12f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.650 2.905 1.235 ;
        RECT 2.245 0.900 2.895 1.225 ;
        RECT 3.300 0.135 3.625 0.72 ;
        RECT 2.580 0.650 3.62 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.755 0.720 1.275 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.720 2.06 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.205 0.740 3.79 0.805 ;
        END
    END c
END oa12f03

MACRO oa12f04
    CLASS CORE ;
    FOREIGN oa12f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.010 0.650 3.4 1.235 ;
        RECT 2.620 0.900 3.4 1.225 ;
        RECT 3.850 0.135 4.24 0.72 ;
        RECT 3.010 0.650 4.245 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.880 0.720 1.465 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.945 0.720 2.4 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.740 0.740 4.455 0.805 ;
        END
    END c
END oa12f04

MACRO oa12f06
    CLASS CORE ;
    FOREIGN oa12f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.655 0.650 4.11 1.235 ;
        RECT 3.180 0.900 4.09 1.225 ;
        RECT 4.675 0.135 5.13 0.72 ;
        RECT 3.655 0.650 5.085 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.070 0.720 1.85 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.365 0.720 2.885 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.540 0.740 5.385 0.805 ;
        END
    END c
END oa12f06

MACRO oa12f08
    CLASS CORE ;
    FOREIGN oa12f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.650 4.82 1.235 ;
        RECT 3.740 0.900 4.845 1.225 ;
        RECT 5.500 0.135 6.02 0.72 ;
        RECT 4.300 0.650 5.99 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.260 0.720 2.17 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.720 3.43 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.340 0.740 6.315 0.805 ;
        END
    END c
END oa12f08

MACRO oa12f10
    CLASS CORE ;
    FOREIGN oa12f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.730 0.650 5.315 1.235 ;
        RECT 4.115 0.900 5.285 1.225 ;
        RECT 6.050 0.135 6.635 0.72 ;
        RECT 4.730 0.650 6.615 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.385 0.720 2.36 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.060 0.720 3.775 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.875 0.740 6.98 0.805 ;
        END
    END c
END oa12f10

MACRO oa12f20
    CLASS CORE ;
    FOREIGN oa12f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.400 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.450 0.650 7.23 1.235 ;
        RECT 5.610 0.900 7.235 1.225 ;
        RECT 8.250 0.135 9.03 0.72 ;
        RECT 6.450 0.650 9.05 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.890 0.720 3.19 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.170 0.720 5.145 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.010 0.740 9.505 0.805 ;
        END
    END c
END oa12f20

MACRO oa12f40
    CLASS CORE ;
    FOREIGN oa12f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.815 0.650 9.855 1.235 ;
        RECT 7.665 0.900 9.875 1.225 ;
        RECT 11.275 0.135 12.315 0.72 ;
        RECT 8.815 0.650 12.325 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.585 0.720 4.405 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.700 0.720 7.0 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.945 0.740 13.025 0.805 ;
        END
    END c
END oa12f40

MACRO oa12f80
    CLASS CORE ;
    FOREIGN oa12f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.255 0.650 13.75 1.235 ;
        RECT 10.660 0.900 13.715 1.225 ;
        RECT 15.675 0.135 17.17 0.72 ;
        RECT 12.255 0.650 17.13 0.715 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.720 6.125 0.785 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.925 0.720 9.745 0.785 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 15.220 0.740 18.08 0.805 ;
        END
    END c
END oa12f80

MACRO oa22s01
    CLASS CORE ;
    FOREIGN oa22s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.210 0.53 0.925 ;
        RECT 0.465 0.870 0.79 0.935 ;
        RECT 0.715 0.870 0.78 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.725 1.34 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.725 1.085 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.635 0.405 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.725 0.83 0.79 ;
        END
    END d
END oa22s01

MACRO oa22s02
    CLASS CORE ;
    FOREIGN oa22s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.180 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.210 1.535 0.925 ;
        RECT 1.275 0.870 2.185 0.935 ;
        RECT 1.970 0.870 2.23 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.145 0.725 3.6 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.445 0.725 2.9 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.580 0.635 1.035 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.750 0.725 2.205 0.79 ;
        END
    END d
END oa22s02

MACRO oa22s03
    CLASS CORE ;
    FOREIGN oa22s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.210 1.945 0.925 ;
        RECT 1.620 0.870 2.79 0.935 ;
        RECT 2.510 0.870 2.835 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.725 4.585 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.725 3.7 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.635 1.32 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.725 2.815 0.79 ;
        END
    END d
END oa22s03

MACRO oa22s04
    CLASS CORE ;
    FOREIGN oa22s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.210 2.18 0.925 ;
        RECT 1.855 0.870 3.22 0.935 ;
        RECT 2.865 0.870 3.19 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.725 5.225 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.725 4.21 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.840 0.635 1.49 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.725 3.195 0.79 ;
        END
    END d
END oa22s04

MACRO oa22s06
    CLASS CORE ;
    FOREIGN oa22s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.220 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.200 0.210 2.59 0.925 ;
        RECT 2.200 0.870 3.825 0.935 ;
        RECT 3.405 0.870 3.795 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.430 0.725 6.21 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.230 0.725 5.01 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.995 0.635 1.775 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.025 0.725 3.805 0.79 ;
        END
    END d
END oa22s06

MACRO oa22s08
    CLASS CORE ;
    FOREIGN oa22s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.550 0.210 3.005 0.925 ;
        RECT 2.550 0.870 4.435 0.935 ;
        RECT 3.940 0.870 4.395 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.290 0.725 7.2 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.895 0.725 5.805 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.155 0.635 2.065 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.500 0.725 4.41 0.79 ;
        END
    END d
END oa22s08

MACRO oa22s10
    CLASS CORE ;
    FOREIGN oa22s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.120 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.210 3.3 0.925 ;
        RECT 2.780 0.870 4.795 0.935 ;
        RECT 4.300 0.870 4.82 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.860 0.725 7.835 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.340 0.725 6.315 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.260 0.635 2.235 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.820 0.725 4.795 0.79 ;
        END
    END d
END oa22s10

MACRO oa22s20
    CLASS CORE ;
    FOREIGN oa22s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.920 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.940 0.210 4.655 0.925 ;
        RECT 3.940 0.870 6.8 0.935 ;
        RECT 6.090 0.870 6.805 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.720 0.725 11.15 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.565 0.725 8.995 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.785 0.635 3.215 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.410 0.725 6.84 0.79 ;
        END
    END d
END oa22s20

MACRO oa22s40
    CLASS CORE ;
    FOREIGN oa22s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.480 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.330 0.210 6.305 0.925 ;
        RECT 5.330 0.870 9.23 0.935 ;
        RECT 8.240 0.870 9.215 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 13.150 0.725 15.035 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.235 0.725 12.12 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.415 0.635 4.3 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.320 0.725 9.205 0.79 ;
        END
    END d
END oa22s40

MACRO oa22s80
    CLASS CORE ;
    FOREIGN oa22s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 24.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.415 0.210 8.78 0.925 ;
        RECT 7.415 0.870 12.875 0.935 ;
        RECT 11.465 0.870 12.83 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 18.295 0.725 20.96 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 14.240 0.725 16.905 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.360 0.635 6.025 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.185 0.725 12.85 0.79 ;
        END
    END d
END oa22s80

MACRO oa22m01
    CLASS CORE ;
    FOREIGN oa22m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.210 0.53 0.925 ;
        RECT 0.465 0.870 0.79 0.935 ;
        RECT 0.715 0.870 0.78 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.725 1.34 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.725 1.085 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.635 0.405 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.725 0.83 0.79 ;
        END
    END d
END oa22m01

MACRO oa22m02
    CLASS CORE ;
    FOREIGN oa22m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.180 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.210 1.535 0.925 ;
        RECT 1.275 0.870 2.185 0.935 ;
        RECT 1.970 0.870 2.23 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.145 0.725 3.6 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.445 0.725 2.9 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.580 0.635 1.035 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.750 0.725 2.205 0.79 ;
        END
    END d
END oa22m02

MACRO oa22m03
    CLASS CORE ;
    FOREIGN oa22m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.210 1.945 0.925 ;
        RECT 1.620 0.870 2.79 0.935 ;
        RECT 2.510 0.870 2.835 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.725 4.585 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.725 3.7 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.635 1.32 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.725 2.815 0.79 ;
        END
    END d
END oa22m03

MACRO oa22m04
    CLASS CORE ;
    FOREIGN oa22m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.210 2.18 0.925 ;
        RECT 1.855 0.870 3.22 0.935 ;
        RECT 2.865 0.870 3.19 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.725 5.225 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.725 4.21 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.840 0.635 1.49 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.725 3.195 0.79 ;
        END
    END d
END oa22m04

MACRO oa22m06
    CLASS CORE ;
    FOREIGN oa22m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.220 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.200 0.210 2.59 0.925 ;
        RECT 2.200 0.870 3.825 0.935 ;
        RECT 3.405 0.870 3.795 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.430 0.725 6.21 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.230 0.725 5.01 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.995 0.635 1.775 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.025 0.725 3.805 0.79 ;
        END
    END d
END oa22m06

MACRO oa22m08
    CLASS CORE ;
    FOREIGN oa22m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.550 0.210 3.005 0.925 ;
        RECT 2.550 0.870 4.435 0.935 ;
        RECT 3.940 0.870 4.395 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.290 0.725 7.2 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.895 0.725 5.805 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.155 0.635 2.065 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.500 0.725 4.41 0.79 ;
        END
    END d
END oa22m08

MACRO oa22m10
    CLASS CORE ;
    FOREIGN oa22m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.120 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.210 3.3 0.925 ;
        RECT 2.780 0.870 4.795 0.935 ;
        RECT 4.300 0.870 4.82 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.860 0.725 7.835 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.340 0.725 6.315 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.260 0.635 2.235 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.820 0.725 4.795 0.79 ;
        END
    END d
END oa22m10

MACRO oa22m20
    CLASS CORE ;
    FOREIGN oa22m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.920 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.940 0.210 4.655 0.925 ;
        RECT 3.940 0.870 6.8 0.935 ;
        RECT 6.090 0.870 6.805 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.720 0.725 11.15 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.565 0.725 8.995 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.785 0.635 3.215 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.410 0.725 6.84 0.79 ;
        END
    END d
END oa22m20

MACRO oa22m40
    CLASS CORE ;
    FOREIGN oa22m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.480 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.330 0.210 6.305 0.925 ;
        RECT 5.330 0.870 9.23 0.935 ;
        RECT 8.240 0.870 9.215 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 13.150 0.725 15.035 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.235 0.725 12.12 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.415 0.635 4.3 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.320 0.725 9.205 0.79 ;
        END
    END d
END oa22m40

MACRO oa22m80
    CLASS CORE ;
    FOREIGN oa22m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 24.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.415 0.210 8.78 0.925 ;
        RECT 7.415 0.870 12.875 0.935 ;
        RECT 11.465 0.870 12.83 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 18.295 0.725 20.96 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 14.240 0.725 16.905 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.360 0.635 6.025 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.185 0.725 12.85 0.79 ;
        END
    END d
END oa22m80

MACRO oa22f01
    CLASS CORE ;
    FOREIGN oa22f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.210 0.53 0.925 ;
        RECT 0.465 0.870 0.79 0.935 ;
        RECT 0.715 0.870 0.78 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.725 1.34 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.725 1.085 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.635 0.405 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.725 0.83 0.79 ;
        END
    END d
END oa22f01

MACRO oa22f02
    CLASS CORE ;
    FOREIGN oa22f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.180 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.210 1.535 0.925 ;
        RECT 1.275 0.870 2.185 0.935 ;
        RECT 1.970 0.870 2.23 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.145 0.725 3.6 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.445 0.725 2.9 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.580 0.635 1.035 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.750 0.725 2.205 0.79 ;
        END
    END d
END oa22f02

MACRO oa22f03
    CLASS CORE ;
    FOREIGN oa22f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.210 1.945 0.925 ;
        RECT 1.620 0.870 2.79 0.935 ;
        RECT 2.510 0.870 2.835 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.725 4.585 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.725 3.7 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.635 1.32 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.725 2.815 0.79 ;
        END
    END d
END oa22f03

MACRO oa22f04
    CLASS CORE ;
    FOREIGN oa22f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.210 2.18 0.925 ;
        RECT 1.855 0.870 3.22 0.935 ;
        RECT 2.865 0.870 3.19 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.725 5.225 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.725 4.21 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.840 0.635 1.49 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.725 3.195 0.79 ;
        END
    END d
END oa22f04

MACRO oa22f06
    CLASS CORE ;
    FOREIGN oa22f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.220 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.200 0.210 2.59 0.925 ;
        RECT 2.200 0.870 3.825 0.935 ;
        RECT 3.405 0.870 3.795 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.430 0.725 6.21 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.230 0.725 5.01 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.995 0.635 1.775 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.025 0.725 3.805 0.79 ;
        END
    END d
END oa22f06

MACRO oa22f08
    CLASS CORE ;
    FOREIGN oa22f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.360 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.550 0.210 3.005 0.925 ;
        RECT 2.550 0.870 4.435 0.935 ;
        RECT 3.940 0.870 4.395 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.290 0.725 7.2 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.895 0.725 5.805 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.155 0.635 2.065 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.500 0.725 4.41 0.79 ;
        END
    END d
END oa22f08

MACRO oa22f10
    CLASS CORE ;
    FOREIGN oa22f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.120 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.210 3.3 0.925 ;
        RECT 2.780 0.870 4.795 0.935 ;
        RECT 4.300 0.870 4.82 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.860 0.725 7.835 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.340 0.725 6.315 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.260 0.635 2.235 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.820 0.725 4.795 0.79 ;
        END
    END d
END oa22f10

MACRO oa22f20
    CLASS CORE ;
    FOREIGN oa22f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.920 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.940 0.210 4.655 0.925 ;
        RECT 3.940 0.870 6.8 0.935 ;
        RECT 6.090 0.870 6.805 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.720 0.725 11.15 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.565 0.725 8.995 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.785 0.635 3.215 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.410 0.725 6.84 0.79 ;
        END
    END d
END oa22f20

MACRO oa22f40
    CLASS CORE ;
    FOREIGN oa22f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.480 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.330 0.210 6.305 0.925 ;
        RECT 5.330 0.870 9.23 0.935 ;
        RECT 8.240 0.870 9.215 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 13.150 0.725 15.035 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.235 0.725 12.12 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.415 0.635 4.3 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.320 0.725 9.205 0.79 ;
        END
    END d
END oa22f40

MACRO oa22f80
    CLASS CORE ;
    FOREIGN oa22f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 24.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 7.415 0.210 8.78 0.925 ;
        RECT 7.415 0.870 12.875 0.935 ;
        RECT 11.465 0.870 12.83 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 18.295 0.725 20.96 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 14.240 0.725 16.905 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.360 0.635 6.025 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 10.185 0.725 12.85 0.79 ;
        END
    END d
END oa22f80

MACRO ms00f80
    CLASS CORE ;
    FOREIGN ms00f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.150 0.150 0.345 1.58 ;
        RECT 0.150 0.635 0.605 0.7 ;
        RECT 0.150 1.140 1.255 1.205 ;
        END
    END o
    PIN ck
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.195 0.990 4.39 1.38 ;
        RECT 4.195 0.990 4.455 1.185 ;
        RECT 1.450 0.640 1.645 0.835 ;
        RECT 1.250 0.780 1.64 0.845 ;
        RECT 1.450 0.640 2.815 0.705 ;
        RECT 2.250 0.640 2.835 0.835 ;
        RECT 3.465 0.705 3.855 0.835 ;
        RECT 2.250 0.790 3.875 0.855 ;
        RECT 3.665 0.705 3.86 1.03 ;
        RECT 3.665 1.015 4.51 1.08 ;
        RECT 4.150 1.015 4.54 1.145 ;
        RECT 4.195 1.290 4.39 1.485 ;
        RECT 6.350 0.775 6.805 0.84 ;
        RECT 6.595 0.775 6.79 1.49 ;
        RECT 4.195 1.470 6.795 1.535 ;
        RECT 4.195 1.315 4.39 1.38 ;
        RECT 4.250 1.110 4.445 1.175 ;
        RECT 4.250 1.015 4.445 1.08 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.965 0.720 7.16 0.785 ;
        END
    END d
END ms00f80

