(* techmap_wrap = "booth" *)
(* techmap_celltype = "$macc" *)
module _70_macc;
endmodule
