module aes_cipher_top (clk,
    rst,
    ld,
    done,
    key,
    text_in,
    text_out);
 input clk;
 input rst;
 input ld;
 output done;
 input [127:0] key;
 input [127:0] text_in;
 output [127:0] text_out;

 FILLCELL_X1 PHY_1 ();
 FILLCELL_X1 PHY_10 ();
 FILLCELL_X1 PHY_100 ();
 FILLCELL_X1 PHY_101 ();
 FILLCELL_X1 PHY_102 ();
 FILLCELL_X1 PHY_103 ();
 FILLCELL_X1 PHY_104 ();
 FILLCELL_X1 PHY_105 ();
 FILLCELL_X1 PHY_106 ();
 FILLCELL_X1 PHY_107 ();
 FILLCELL_X1 PHY_108 ();
 FILLCELL_X1 PHY_109 ();
 FILLCELL_X1 PHY_11 ();
 FILLCELL_X1 PHY_110 ();
 FILLCELL_X1 PHY_111 ();
 FILLCELL_X1 PHY_112 ();
 FILLCELL_X1 PHY_113 ();
 FILLCELL_X1 PHY_114 ();
 FILLCELL_X1 PHY_115 ();
 FILLCELL_X1 PHY_116 ();
 FILLCELL_X1 PHY_117 ();
 FILLCELL_X1 PHY_118 ();
 FILLCELL_X1 PHY_119 ();
 FILLCELL_X1 PHY_12 ();
 FILLCELL_X1 PHY_120 ();
 FILLCELL_X1 PHY_121 ();
 FILLCELL_X1 PHY_122 ();
 FILLCELL_X1 PHY_123 ();
 FILLCELL_X1 PHY_124 ();
 FILLCELL_X1 PHY_125 ();
 FILLCELL_X1 PHY_126 ();
 FILLCELL_X1 PHY_127 ();
 FILLCELL_X1 PHY_128 ();
 FILLCELL_X1 PHY_129 ();
 FILLCELL_X1 PHY_13 ();
 FILLCELL_X1 PHY_130 ();
 FILLCELL_X1 PHY_131 ();
 FILLCELL_X1 PHY_132 ();
 FILLCELL_X1 PHY_133 ();
 FILLCELL_X1 PHY_134 ();
 FILLCELL_X1 PHY_135 ();
 FILLCELL_X1 PHY_136 ();
 FILLCELL_X1 PHY_137 ();
 FILLCELL_X1 PHY_138 ();
 FILLCELL_X1 PHY_139 ();
 FILLCELL_X1 PHY_14 ();
 FILLCELL_X1 PHY_140 ();
 FILLCELL_X1 PHY_141 ();
 FILLCELL_X1 PHY_142 ();
 FILLCELL_X1 PHY_143 ();
 FILLCELL_X1 PHY_144 ();
 FILLCELL_X1 PHY_145 ();
 FILLCELL_X1 PHY_146 ();
 FILLCELL_X1 PHY_147 ();
 FILLCELL_X1 PHY_148 ();
 FILLCELL_X1 PHY_149 ();
 FILLCELL_X1 PHY_15 ();
 FILLCELL_X1 PHY_150 ();
 FILLCELL_X1 PHY_151 ();
 FILLCELL_X1 PHY_152 ();
 FILLCELL_X1 PHY_153 ();
 FILLCELL_X1 PHY_154 ();
 FILLCELL_X1 PHY_155 ();
 FILLCELL_X1 PHY_156 ();
 FILLCELL_X1 PHY_157 ();
 FILLCELL_X1 PHY_158 ();
 FILLCELL_X1 PHY_159 ();
 FILLCELL_X1 PHY_16 ();
 FILLCELL_X1 PHY_160 ();
 FILLCELL_X1 PHY_161 ();
 FILLCELL_X1 PHY_162 ();
 FILLCELL_X1 PHY_163 ();
 FILLCELL_X1 PHY_164 ();
 FILLCELL_X1 PHY_165 ();
 FILLCELL_X1 PHY_166 ();
 FILLCELL_X1 PHY_167 ();
 FILLCELL_X1 PHY_168 ();
 FILLCELL_X1 PHY_169 ();
 FILLCELL_X1 PHY_17 ();
 FILLCELL_X1 PHY_170 ();
 FILLCELL_X1 PHY_171 ();
 FILLCELL_X1 PHY_172 ();
 FILLCELL_X1 PHY_173 ();
 FILLCELL_X1 PHY_174 ();
 FILLCELL_X1 PHY_175 ();
 FILLCELL_X1 PHY_176 ();
 FILLCELL_X1 PHY_177 ();
 FILLCELL_X1 PHY_178 ();
 FILLCELL_X1 PHY_179 ();
 FILLCELL_X1 PHY_18 ();
 FILLCELL_X1 PHY_180 ();
 FILLCELL_X1 PHY_181 ();
 FILLCELL_X1 PHY_182 ();
 FILLCELL_X1 PHY_183 ();
 FILLCELL_X1 PHY_184 ();
 FILLCELL_X1 PHY_185 ();
 FILLCELL_X1 PHY_186 ();
 FILLCELL_X1 PHY_187 ();
 FILLCELL_X1 PHY_188 ();
 FILLCELL_X1 PHY_189 ();
 FILLCELL_X1 PHY_19 ();
 FILLCELL_X1 PHY_190 ();
 FILLCELL_X1 PHY_191 ();
 FILLCELL_X1 PHY_192 ();
 FILLCELL_X1 PHY_193 ();
 FILLCELL_X1 PHY_194 ();
 FILLCELL_X1 PHY_195 ();
 FILLCELL_X1 PHY_196 ();
 FILLCELL_X1 PHY_197 ();
 FILLCELL_X1 PHY_198 ();
 FILLCELL_X1 PHY_199 ();
 FILLCELL_X1 PHY_2 ();
 FILLCELL_X1 PHY_20 ();
 FILLCELL_X1 PHY_200 ();
 FILLCELL_X1 PHY_201 ();
 FILLCELL_X1 PHY_202 ();
 FILLCELL_X1 PHY_203 ();
 FILLCELL_X1 PHY_204 ();
 FILLCELL_X1 PHY_205 ();
 FILLCELL_X1 PHY_206 ();
 FILLCELL_X1 PHY_207 ();
 FILLCELL_X1 PHY_208 ();
 FILLCELL_X1 PHY_209 ();
 FILLCELL_X1 PHY_21 ();
 FILLCELL_X1 PHY_210 ();
 FILLCELL_X1 PHY_211 ();
 FILLCELL_X1 PHY_212 ();
 FILLCELL_X1 PHY_213 ();
 FILLCELL_X1 PHY_214 ();
 FILLCELL_X1 PHY_215 ();
 FILLCELL_X1 PHY_216 ();
 FILLCELL_X1 PHY_217 ();
 FILLCELL_X1 PHY_218 ();
 FILLCELL_X1 PHY_219 ();
 FILLCELL_X1 PHY_22 ();
 FILLCELL_X1 PHY_220 ();
 FILLCELL_X1 PHY_221 ();
 FILLCELL_X1 PHY_222 ();
 FILLCELL_X1 PHY_223 ();
 FILLCELL_X1 PHY_224 ();
 FILLCELL_X1 PHY_225 ();
 FILLCELL_X1 PHY_226 ();
 FILLCELL_X1 PHY_227 ();
 FILLCELL_X1 PHY_228 ();
 FILLCELL_X1 PHY_229 ();
 FILLCELL_X1 PHY_23 ();
 FILLCELL_X1 PHY_230 ();
 FILLCELL_X1 PHY_231 ();
 FILLCELL_X1 PHY_232 ();
 FILLCELL_X1 PHY_233 ();
 FILLCELL_X1 PHY_234 ();
 FILLCELL_X1 PHY_235 ();
 FILLCELL_X1 PHY_236 ();
 FILLCELL_X1 PHY_237 ();
 FILLCELL_X1 PHY_238 ();
 FILLCELL_X1 PHY_239 ();
 FILLCELL_X1 PHY_24 ();
 FILLCELL_X1 PHY_240 ();
 FILLCELL_X1 PHY_241 ();
 FILLCELL_X1 PHY_242 ();
 FILLCELL_X1 PHY_243 ();
 FILLCELL_X1 PHY_244 ();
 FILLCELL_X1 PHY_245 ();
 FILLCELL_X1 PHY_246 ();
 FILLCELL_X1 PHY_247 ();
 FILLCELL_X1 PHY_248 ();
 FILLCELL_X1 PHY_249 ();
 FILLCELL_X1 PHY_25 ();
 FILLCELL_X1 PHY_250 ();
 FILLCELL_X1 PHY_251 ();
 FILLCELL_X1 PHY_252 ();
 FILLCELL_X1 PHY_253 ();
 FILLCELL_X1 PHY_254 ();
 FILLCELL_X1 PHY_255 ();
 FILLCELL_X1 PHY_256 ();
 FILLCELL_X1 PHY_257 ();
 FILLCELL_X1 PHY_258 ();
 FILLCELL_X1 PHY_259 ();
 FILLCELL_X1 PHY_26 ();
 FILLCELL_X1 PHY_260 ();
 FILLCELL_X1 PHY_261 ();
 FILLCELL_X1 PHY_262 ();
 FILLCELL_X1 PHY_263 ();
 FILLCELL_X1 PHY_264 ();
 FILLCELL_X1 PHY_265 ();
 FILLCELL_X1 PHY_266 ();
 FILLCELL_X1 PHY_267 ();
 FILLCELL_X1 PHY_268 ();
 FILLCELL_X1 PHY_269 ();
 FILLCELL_X1 PHY_27 ();
 FILLCELL_X1 PHY_270 ();
 FILLCELL_X1 PHY_271 ();
 FILLCELL_X1 PHY_272 ();
 FILLCELL_X1 PHY_273 ();
 FILLCELL_X1 PHY_274 ();
 FILLCELL_X1 PHY_275 ();
 FILLCELL_X1 PHY_276 ();
 FILLCELL_X1 PHY_277 ();
 FILLCELL_X1 PHY_278 ();
 FILLCELL_X1 PHY_279 ();
 FILLCELL_X1 PHY_28 ();
 FILLCELL_X1 PHY_280 ();
 FILLCELL_X1 PHY_281 ();
 FILLCELL_X1 PHY_282 ();
 FILLCELL_X1 PHY_283 ();
 FILLCELL_X1 PHY_284 ();
 FILLCELL_X1 PHY_285 ();
 FILLCELL_X1 PHY_286 ();
 FILLCELL_X1 PHY_287 ();
 FILLCELL_X1 PHY_288 ();
 FILLCELL_X1 PHY_289 ();
 FILLCELL_X1 PHY_29 ();
 FILLCELL_X1 PHY_290 ();
 FILLCELL_X1 PHY_291 ();
 FILLCELL_X1 PHY_292 ();
 FILLCELL_X1 PHY_293 ();
 FILLCELL_X1 PHY_294 ();
 FILLCELL_X1 PHY_295 ();
 FILLCELL_X1 PHY_296 ();
 FILLCELL_X1 PHY_297 ();
 FILLCELL_X1 PHY_298 ();
 FILLCELL_X1 PHY_299 ();
 FILLCELL_X1 PHY_3 ();
 FILLCELL_X1 PHY_30 ();
 FILLCELL_X1 PHY_300 ();
 FILLCELL_X1 PHY_301 ();
 FILLCELL_X1 PHY_302 ();
 FILLCELL_X1 PHY_303 ();
 FILLCELL_X1 PHY_304 ();
 FILLCELL_X1 PHY_305 ();
 FILLCELL_X1 PHY_306 ();
 FILLCELL_X1 PHY_307 ();
 FILLCELL_X1 PHY_308 ();
 FILLCELL_X1 PHY_309 ();
 FILLCELL_X1 PHY_31 ();
 FILLCELL_X1 PHY_310 ();
 FILLCELL_X1 PHY_311 ();
 FILLCELL_X1 PHY_312 ();
 FILLCELL_X1 PHY_313 ();
 FILLCELL_X1 PHY_314 ();
 FILLCELL_X1 PHY_315 ();
 FILLCELL_X1 PHY_316 ();
 FILLCELL_X1 PHY_317 ();
 FILLCELL_X1 PHY_318 ();
 FILLCELL_X1 PHY_319 ();
 FILLCELL_X1 PHY_32 ();
 FILLCELL_X1 PHY_320 ();
 FILLCELL_X1 PHY_321 ();
 FILLCELL_X1 PHY_322 ();
 FILLCELL_X1 PHY_323 ();
 FILLCELL_X1 PHY_324 ();
 FILLCELL_X1 PHY_325 ();
 FILLCELL_X1 PHY_326 ();
 FILLCELL_X1 PHY_327 ();
 FILLCELL_X1 PHY_328 ();
 FILLCELL_X1 PHY_329 ();
 FILLCELL_X1 PHY_33 ();
 FILLCELL_X1 PHY_330 ();
 FILLCELL_X1 PHY_331 ();
 FILLCELL_X1 PHY_332 ();
 FILLCELL_X1 PHY_333 ();
 FILLCELL_X1 PHY_334 ();
 FILLCELL_X1 PHY_335 ();
 FILLCELL_X1 PHY_336 ();
 FILLCELL_X1 PHY_337 ();
 FILLCELL_X1 PHY_338 ();
 FILLCELL_X1 PHY_339 ();
 FILLCELL_X1 PHY_34 ();
 FILLCELL_X1 PHY_340 ();
 FILLCELL_X1 PHY_341 ();
 FILLCELL_X1 PHY_342 ();
 FILLCELL_X1 PHY_343 ();
 FILLCELL_X1 PHY_344 ();
 FILLCELL_X1 PHY_345 ();
 FILLCELL_X1 PHY_346 ();
 FILLCELL_X1 PHY_347 ();
 FILLCELL_X1 PHY_348 ();
 FILLCELL_X1 PHY_349 ();
 FILLCELL_X1 PHY_35 ();
 FILLCELL_X1 PHY_350 ();
 FILLCELL_X1 PHY_351 ();
 FILLCELL_X1 PHY_352 ();
 FILLCELL_X1 PHY_353 ();
 FILLCELL_X1 PHY_354 ();
 FILLCELL_X1 PHY_355 ();
 FILLCELL_X1 PHY_356 ();
 FILLCELL_X1 PHY_357 ();
 FILLCELL_X1 PHY_358 ();
 FILLCELL_X1 PHY_359 ();
 FILLCELL_X1 PHY_36 ();
 FILLCELL_X1 PHY_360 ();
 FILLCELL_X1 PHY_361 ();
 FILLCELL_X1 PHY_362 ();
 FILLCELL_X1 PHY_363 ();
 FILLCELL_X1 PHY_364 ();
 FILLCELL_X1 PHY_365 ();
 FILLCELL_X1 PHY_366 ();
 FILLCELL_X1 PHY_367 ();
 FILLCELL_X1 PHY_368 ();
 FILLCELL_X1 PHY_369 ();
 FILLCELL_X1 PHY_37 ();
 FILLCELL_X1 PHY_370 ();
 FILLCELL_X1 PHY_371 ();
 FILLCELL_X1 PHY_372 ();
 FILLCELL_X1 PHY_373 ();
 FILLCELL_X1 PHY_374 ();
 FILLCELL_X1 PHY_375 ();
 FILLCELL_X1 PHY_376 ();
 FILLCELL_X1 PHY_377 ();
 FILLCELL_X1 PHY_378 ();
 FILLCELL_X1 PHY_379 ();
 FILLCELL_X1 PHY_38 ();
 FILLCELL_X1 PHY_380 ();
 FILLCELL_X1 PHY_381 ();
 FILLCELL_X1 PHY_382 ();
 FILLCELL_X1 PHY_383 ();
 FILLCELL_X1 PHY_384 ();
 FILLCELL_X1 PHY_385 ();
 FILLCELL_X1 PHY_386 ();
 FILLCELL_X1 PHY_387 ();
 FILLCELL_X1 PHY_388 ();
 FILLCELL_X1 PHY_389 ();
 FILLCELL_X1 PHY_39 ();
 FILLCELL_X1 PHY_390 ();
 FILLCELL_X1 PHY_391 ();
 FILLCELL_X1 PHY_392 ();
 FILLCELL_X1 PHY_393 ();
 FILLCELL_X1 PHY_394 ();
 FILLCELL_X1 PHY_395 ();
 FILLCELL_X1 PHY_396 ();
 FILLCELL_X1 PHY_397 ();
 FILLCELL_X1 PHY_398 ();
 FILLCELL_X1 PHY_399 ();
 FILLCELL_X1 PHY_4 ();
 FILLCELL_X1 PHY_40 ();
 FILLCELL_X1 PHY_400 ();
 FILLCELL_X1 PHY_401 ();
 FILLCELL_X1 PHY_402 ();
 FILLCELL_X1 PHY_403 ();
 FILLCELL_X1 PHY_404 ();
 FILLCELL_X1 PHY_405 ();
 FILLCELL_X1 PHY_406 ();
 FILLCELL_X1 PHY_407 ();
 FILLCELL_X1 PHY_408 ();
 FILLCELL_X1 PHY_409 ();
 FILLCELL_X1 PHY_41 ();
 FILLCELL_X1 PHY_410 ();
 FILLCELL_X1 PHY_411 ();
 FILLCELL_X1 PHY_412 ();
 FILLCELL_X1 PHY_413 ();
 FILLCELL_X1 PHY_414 ();
 FILLCELL_X1 PHY_415 ();
 FILLCELL_X1 PHY_416 ();
 FILLCELL_X1 PHY_417 ();
 FILLCELL_X1 PHY_418 ();
 FILLCELL_X1 PHY_419 ();
 FILLCELL_X1 PHY_42 ();
 FILLCELL_X1 PHY_420 ();
 FILLCELL_X1 PHY_421 ();
 FILLCELL_X1 PHY_422 ();
 FILLCELL_X1 PHY_423 ();
 FILLCELL_X1 PHY_424 ();
 FILLCELL_X1 PHY_425 ();
 FILLCELL_X1 PHY_426 ();
 FILLCELL_X1 PHY_427 ();
 FILLCELL_X1 PHY_428 ();
 FILLCELL_X1 PHY_429 ();
 FILLCELL_X1 PHY_43 ();
 FILLCELL_X1 PHY_430 ();
 FILLCELL_X1 PHY_431 ();
 FILLCELL_X1 PHY_432 ();
 FILLCELL_X1 PHY_433 ();
 FILLCELL_X1 PHY_434 ();
 FILLCELL_X1 PHY_435 ();
 FILLCELL_X1 PHY_436 ();
 FILLCELL_X1 PHY_437 ();
 FILLCELL_X1 PHY_438 ();
 FILLCELL_X1 PHY_439 ();
 FILLCELL_X1 PHY_44 ();
 FILLCELL_X1 PHY_440 ();
 FILLCELL_X1 PHY_441 ();
 FILLCELL_X1 PHY_442 ();
 FILLCELL_X1 PHY_443 ();
 FILLCELL_X1 PHY_444 ();
 FILLCELL_X1 PHY_445 ();
 FILLCELL_X1 PHY_446 ();
 FILLCELL_X1 PHY_447 ();
 FILLCELL_X1 PHY_448 ();
 FILLCELL_X1 PHY_449 ();
 FILLCELL_X1 PHY_45 ();
 FILLCELL_X1 PHY_450 ();
 FILLCELL_X1 PHY_451 ();
 FILLCELL_X1 PHY_452 ();
 FILLCELL_X1 PHY_453 ();
 FILLCELL_X1 PHY_454 ();
 FILLCELL_X1 PHY_455 ();
 FILLCELL_X1 PHY_456 ();
 FILLCELL_X1 PHY_457 ();
 FILLCELL_X1 PHY_458 ();
 FILLCELL_X1 PHY_459 ();
 FILLCELL_X1 PHY_46 ();
 FILLCELL_X1 PHY_460 ();
 FILLCELL_X1 PHY_461 ();
 FILLCELL_X1 PHY_462 ();
 FILLCELL_X1 PHY_463 ();
 FILLCELL_X1 PHY_464 ();
 FILLCELL_X1 PHY_465 ();
 FILLCELL_X1 PHY_466 ();
 FILLCELL_X1 PHY_467 ();
 FILLCELL_X1 PHY_468 ();
 FILLCELL_X1 PHY_469 ();
 FILLCELL_X1 PHY_47 ();
 FILLCELL_X1 PHY_470 ();
 FILLCELL_X1 PHY_471 ();
 FILLCELL_X1 PHY_472 ();
 FILLCELL_X1 PHY_473 ();
 FILLCELL_X1 PHY_474 ();
 FILLCELL_X1 PHY_475 ();
 FILLCELL_X1 PHY_476 ();
 FILLCELL_X1 PHY_477 ();
 FILLCELL_X1 PHY_478 ();
 FILLCELL_X1 PHY_479 ();
 FILLCELL_X1 PHY_48 ();
 FILLCELL_X1 PHY_480 ();
 FILLCELL_X1 PHY_481 ();
 FILLCELL_X1 PHY_482 ();
 FILLCELL_X1 PHY_483 ();
 FILLCELL_X1 PHY_484 ();
 FILLCELL_X1 PHY_485 ();
 FILLCELL_X1 PHY_486 ();
 FILLCELL_X1 PHY_487 ();
 FILLCELL_X1 PHY_488 ();
 FILLCELL_X1 PHY_489 ();
 FILLCELL_X1 PHY_49 ();
 FILLCELL_X1 PHY_490 ();
 FILLCELL_X1 PHY_491 ();
 FILLCELL_X1 PHY_492 ();
 FILLCELL_X1 PHY_493 ();
 FILLCELL_X1 PHY_494 ();
 FILLCELL_X1 PHY_495 ();
 FILLCELL_X1 PHY_496 ();
 FILLCELL_X1 PHY_497 ();
 FILLCELL_X1 PHY_498 ();
 FILLCELL_X1 PHY_499 ();
 FILLCELL_X1 PHY_5 ();
 FILLCELL_X1 PHY_50 ();
 FILLCELL_X1 PHY_500 ();
 FILLCELL_X1 PHY_501 ();
 FILLCELL_X1 PHY_502 ();
 FILLCELL_X1 PHY_503 ();
 FILLCELL_X1 PHY_504 ();
 FILLCELL_X1 PHY_505 ();
 FILLCELL_X1 PHY_506 ();
 FILLCELL_X1 PHY_507 ();
 FILLCELL_X1 PHY_508 ();
 FILLCELL_X1 PHY_509 ();
 FILLCELL_X1 PHY_51 ();
 FILLCELL_X1 PHY_510 ();
 FILLCELL_X1 PHY_511 ();
 FILLCELL_X1 PHY_512 ();
 FILLCELL_X1 PHY_513 ();
 FILLCELL_X1 PHY_514 ();
 FILLCELL_X1 PHY_515 ();
 FILLCELL_X1 PHY_516 ();
 FILLCELL_X1 PHY_517 ();
 FILLCELL_X1 PHY_518 ();
 FILLCELL_X1 PHY_519 ();
 FILLCELL_X1 PHY_52 ();
 FILLCELL_X1 PHY_520 ();
 FILLCELL_X1 PHY_521 ();
 FILLCELL_X1 PHY_522 ();
 FILLCELL_X1 PHY_523 ();
 FILLCELL_X1 PHY_524 ();
 FILLCELL_X1 PHY_525 ();
 FILLCELL_X1 PHY_526 ();
 FILLCELL_X1 PHY_527 ();
 FILLCELL_X1 PHY_528 ();
 FILLCELL_X1 PHY_529 ();
 FILLCELL_X1 PHY_53 ();
 FILLCELL_X1 PHY_530 ();
 FILLCELL_X1 PHY_531 ();
 FILLCELL_X1 PHY_532 ();
 FILLCELL_X1 PHY_533 ();
 FILLCELL_X1 PHY_534 ();
 FILLCELL_X1 PHY_535 ();
 FILLCELL_X1 PHY_536 ();
 FILLCELL_X1 PHY_537 ();
 FILLCELL_X1 PHY_538 ();
 FILLCELL_X1 PHY_539 ();
 FILLCELL_X1 PHY_54 ();
 FILLCELL_X1 PHY_540 ();
 FILLCELL_X1 PHY_541 ();
 FILLCELL_X1 PHY_542 ();
 FILLCELL_X1 PHY_543 ();
 FILLCELL_X1 PHY_544 ();
 FILLCELL_X1 PHY_545 ();
 FILLCELL_X1 PHY_546 ();
 FILLCELL_X1 PHY_547 ();
 FILLCELL_X1 PHY_548 ();
 FILLCELL_X1 PHY_549 ();
 FILLCELL_X1 PHY_55 ();
 FILLCELL_X1 PHY_550 ();
 FILLCELL_X1 PHY_551 ();
 FILLCELL_X1 PHY_552 ();
 FILLCELL_X1 PHY_553 ();
 FILLCELL_X1 PHY_554 ();
 FILLCELL_X1 PHY_555 ();
 FILLCELL_X1 PHY_556 ();
 FILLCELL_X1 PHY_557 ();
 FILLCELL_X1 PHY_558 ();
 FILLCELL_X1 PHY_559 ();
 FILLCELL_X1 PHY_56 ();
 FILLCELL_X1 PHY_560 ();
 FILLCELL_X1 PHY_561 ();
 FILLCELL_X1 PHY_562 ();
 FILLCELL_X1 PHY_563 ();
 FILLCELL_X1 PHY_564 ();
 FILLCELL_X1 PHY_565 ();
 FILLCELL_X1 PHY_566 ();
 FILLCELL_X1 PHY_567 ();
 FILLCELL_X1 PHY_568 ();
 FILLCELL_X1 PHY_569 ();
 FILLCELL_X1 PHY_57 ();
 FILLCELL_X1 PHY_570 ();
 FILLCELL_X1 PHY_571 ();
 FILLCELL_X1 PHY_572 ();
 FILLCELL_X1 PHY_573 ();
 FILLCELL_X1 PHY_574 ();
 FILLCELL_X1 PHY_575 ();
 FILLCELL_X1 PHY_576 ();
 FILLCELL_X1 PHY_577 ();
 FILLCELL_X1 PHY_578 ();
 FILLCELL_X1 PHY_579 ();
 FILLCELL_X1 PHY_58 ();
 FILLCELL_X1 PHY_580 ();
 FILLCELL_X1 PHY_581 ();
 FILLCELL_X1 PHY_582 ();
 FILLCELL_X1 PHY_583 ();
 FILLCELL_X1 PHY_584 ();
 FILLCELL_X1 PHY_585 ();
 FILLCELL_X1 PHY_586 ();
 FILLCELL_X1 PHY_587 ();
 FILLCELL_X1 PHY_588 ();
 FILLCELL_X1 PHY_589 ();
 FILLCELL_X1 PHY_59 ();
 FILLCELL_X1 PHY_590 ();
 FILLCELL_X1 PHY_591 ();
 FILLCELL_X1 PHY_592 ();
 FILLCELL_X1 PHY_593 ();
 FILLCELL_X1 PHY_594 ();
 FILLCELL_X1 PHY_595 ();
 FILLCELL_X1 PHY_596 ();
 FILLCELL_X1 PHY_597 ();
 FILLCELL_X1 PHY_598 ();
 FILLCELL_X1 PHY_599 ();
 FILLCELL_X1 PHY_6 ();
 FILLCELL_X1 PHY_60 ();
 FILLCELL_X1 PHY_600 ();
 FILLCELL_X1 PHY_601 ();
 FILLCELL_X1 PHY_602 ();
 FILLCELL_X1 PHY_603 ();
 FILLCELL_X1 PHY_604 ();
 FILLCELL_X1 PHY_605 ();
 FILLCELL_X1 PHY_606 ();
 FILLCELL_X1 PHY_607 ();
 FILLCELL_X1 PHY_608 ();
 FILLCELL_X1 PHY_609 ();
 FILLCELL_X1 PHY_61 ();
 FILLCELL_X1 PHY_610 ();
 FILLCELL_X1 PHY_611 ();
 FILLCELL_X1 PHY_612 ();
 FILLCELL_X1 PHY_613 ();
 FILLCELL_X1 PHY_614 ();
 FILLCELL_X1 PHY_615 ();
 FILLCELL_X1 PHY_616 ();
 FILLCELL_X1 PHY_617 ();
 FILLCELL_X1 PHY_618 ();
 FILLCELL_X1 PHY_619 ();
 FILLCELL_X1 PHY_62 ();
 FILLCELL_X1 PHY_620 ();
 FILLCELL_X1 PHY_621 ();
 FILLCELL_X1 PHY_622 ();
 FILLCELL_X1 PHY_623 ();
 FILLCELL_X1 PHY_624 ();
 FILLCELL_X1 PHY_625 ();
 FILLCELL_X1 PHY_626 ();
 FILLCELL_X1 PHY_627 ();
 FILLCELL_X1 PHY_628 ();
 FILLCELL_X1 PHY_629 ();
 FILLCELL_X1 PHY_63 ();
 FILLCELL_X1 PHY_630 ();
 FILLCELL_X1 PHY_631 ();
 FILLCELL_X1 PHY_632 ();
 FILLCELL_X1 PHY_633 ();
 FILLCELL_X1 PHY_634 ();
 FILLCELL_X1 PHY_635 ();
 FILLCELL_X1 PHY_636 ();
 FILLCELL_X1 PHY_637 ();
 FILLCELL_X1 PHY_638 ();
 FILLCELL_X1 PHY_639 ();
 FILLCELL_X1 PHY_64 ();
 FILLCELL_X1 PHY_640 ();
 FILLCELL_X1 PHY_641 ();
 FILLCELL_X1 PHY_642 ();
 FILLCELL_X1 PHY_643 ();
 FILLCELL_X1 PHY_644 ();
 FILLCELL_X1 PHY_645 ();
 FILLCELL_X1 PHY_646 ();
 FILLCELL_X1 PHY_647 ();
 FILLCELL_X1 PHY_648 ();
 FILLCELL_X1 PHY_649 ();
 FILLCELL_X1 PHY_65 ();
 FILLCELL_X1 PHY_650 ();
 FILLCELL_X1 PHY_651 ();
 FILLCELL_X1 PHY_652 ();
 FILLCELL_X1 PHY_653 ();
 FILLCELL_X1 PHY_654 ();
 FILLCELL_X1 PHY_655 ();
 FILLCELL_X1 PHY_656 ();
 FILLCELL_X1 PHY_657 ();
 FILLCELL_X1 PHY_658 ();
 FILLCELL_X1 PHY_659 ();
 FILLCELL_X1 PHY_66 ();
 FILLCELL_X1 PHY_660 ();
 FILLCELL_X1 PHY_661 ();
 FILLCELL_X1 PHY_662 ();
 FILLCELL_X1 PHY_663 ();
 FILLCELL_X1 PHY_664 ();
 FILLCELL_X1 PHY_665 ();
 FILLCELL_X1 PHY_666 ();
 FILLCELL_X1 PHY_667 ();
 FILLCELL_X1 PHY_668 ();
 FILLCELL_X1 PHY_669 ();
 FILLCELL_X1 PHY_67 ();
 FILLCELL_X1 PHY_670 ();
 FILLCELL_X1 PHY_671 ();
 FILLCELL_X1 PHY_672 ();
 FILLCELL_X1 PHY_673 ();
 FILLCELL_X1 PHY_674 ();
 FILLCELL_X1 PHY_675 ();
 FILLCELL_X1 PHY_676 ();
 FILLCELL_X1 PHY_677 ();
 FILLCELL_X1 PHY_678 ();
 FILLCELL_X1 PHY_679 ();
 FILLCELL_X1 PHY_68 ();
 FILLCELL_X1 PHY_680 ();
 FILLCELL_X1 PHY_681 ();
 FILLCELL_X1 PHY_682 ();
 FILLCELL_X1 PHY_683 ();
 FILLCELL_X1 PHY_684 ();
 FILLCELL_X1 PHY_685 ();
 FILLCELL_X1 PHY_686 ();
 FILLCELL_X1 PHY_687 ();
 FILLCELL_X1 PHY_688 ();
 FILLCELL_X1 PHY_689 ();
 FILLCELL_X1 PHY_69 ();
 FILLCELL_X1 PHY_690 ();
 FILLCELL_X1 PHY_691 ();
 FILLCELL_X1 PHY_692 ();
 FILLCELL_X1 PHY_693 ();
 FILLCELL_X1 PHY_694 ();
 FILLCELL_X1 PHY_695 ();
 FILLCELL_X1 PHY_696 ();
 FILLCELL_X1 PHY_697 ();
 FILLCELL_X1 PHY_698 ();
 FILLCELL_X1 PHY_699 ();
 FILLCELL_X1 PHY_7 ();
 FILLCELL_X1 PHY_70 ();
 FILLCELL_X1 PHY_700 ();
 FILLCELL_X1 PHY_701 ();
 FILLCELL_X1 PHY_702 ();
 FILLCELL_X1 PHY_703 ();
 FILLCELL_X1 PHY_704 ();
 FILLCELL_X1 PHY_705 ();
 FILLCELL_X1 PHY_706 ();
 FILLCELL_X1 PHY_707 ();
 FILLCELL_X1 PHY_708 ();
 FILLCELL_X1 PHY_709 ();
 FILLCELL_X1 PHY_71 ();
 FILLCELL_X1 PHY_710 ();
 FILLCELL_X1 PHY_711 ();
 FILLCELL_X1 PHY_712 ();
 FILLCELL_X1 PHY_713 ();
 FILLCELL_X1 PHY_714 ();
 FILLCELL_X1 PHY_715 ();
 FILLCELL_X1 PHY_716 ();
 FILLCELL_X1 PHY_717 ();
 FILLCELL_X1 PHY_718 ();
 FILLCELL_X1 PHY_719 ();
 FILLCELL_X1 PHY_72 ();
 FILLCELL_X1 PHY_720 ();
 FILLCELL_X1 PHY_721 ();
 FILLCELL_X1 PHY_722 ();
 FILLCELL_X1 PHY_723 ();
 FILLCELL_X1 PHY_724 ();
 FILLCELL_X1 PHY_725 ();
 FILLCELL_X1 PHY_726 ();
 FILLCELL_X1 PHY_727 ();
 FILLCELL_X1 PHY_728 ();
 FILLCELL_X1 PHY_729 ();
 FILLCELL_X1 PHY_73 ();
 FILLCELL_X1 PHY_730 ();
 FILLCELL_X1 PHY_731 ();
 FILLCELL_X1 PHY_732 ();
 FILLCELL_X1 PHY_733 ();
 FILLCELL_X1 PHY_734 ();
 FILLCELL_X1 PHY_735 ();
 FILLCELL_X1 PHY_736 ();
 FILLCELL_X1 PHY_737 ();
 FILLCELL_X1 PHY_738 ();
 FILLCELL_X1 PHY_739 ();
 FILLCELL_X1 PHY_74 ();
 FILLCELL_X1 PHY_740 ();
 FILLCELL_X1 PHY_741 ();
 FILLCELL_X1 PHY_742 ();
 FILLCELL_X1 PHY_743 ();
 FILLCELL_X1 PHY_744 ();
 FILLCELL_X1 PHY_745 ();
 FILLCELL_X1 PHY_746 ();
 FILLCELL_X1 PHY_747 ();
 FILLCELL_X1 PHY_748 ();
 FILLCELL_X1 PHY_749 ();
 FILLCELL_X1 PHY_75 ();
 FILLCELL_X1 PHY_750 ();
 FILLCELL_X1 PHY_751 ();
 FILLCELL_X1 PHY_752 ();
 FILLCELL_X1 PHY_753 ();
 FILLCELL_X1 PHY_754 ();
 FILLCELL_X1 PHY_755 ();
 FILLCELL_X1 PHY_756 ();
 FILLCELL_X1 PHY_757 ();
 FILLCELL_X1 PHY_758 ();
 FILLCELL_X1 PHY_759 ();
 FILLCELL_X1 PHY_76 ();
 FILLCELL_X1 PHY_760 ();
 FILLCELL_X1 PHY_761 ();
 FILLCELL_X1 PHY_762 ();
 FILLCELL_X1 PHY_763 ();
 FILLCELL_X1 PHY_764 ();
 FILLCELL_X1 PHY_765 ();
 FILLCELL_X1 PHY_766 ();
 FILLCELL_X1 PHY_767 ();
 FILLCELL_X1 PHY_768 ();
 FILLCELL_X1 PHY_769 ();
 FILLCELL_X1 PHY_77 ();
 FILLCELL_X1 PHY_770 ();
 FILLCELL_X1 PHY_771 ();
 FILLCELL_X1 PHY_772 ();
 FILLCELL_X1 PHY_773 ();
 FILLCELL_X1 PHY_774 ();
 FILLCELL_X1 PHY_775 ();
 FILLCELL_X1 PHY_776 ();
 FILLCELL_X1 PHY_777 ();
 FILLCELL_X1 PHY_778 ();
 FILLCELL_X1 PHY_779 ();
 FILLCELL_X1 PHY_78 ();
 FILLCELL_X1 PHY_780 ();
 FILLCELL_X1 PHY_781 ();
 FILLCELL_X1 PHY_782 ();
 FILLCELL_X1 PHY_783 ();
 FILLCELL_X1 PHY_784 ();
 FILLCELL_X1 PHY_785 ();
 FILLCELL_X1 PHY_786 ();
 FILLCELL_X1 PHY_787 ();
 FILLCELL_X1 PHY_788 ();
 FILLCELL_X1 PHY_789 ();
 FILLCELL_X1 PHY_79 ();
 FILLCELL_X1 PHY_790 ();
 FILLCELL_X1 PHY_791 ();
 FILLCELL_X1 PHY_792 ();
 FILLCELL_X1 PHY_793 ();
 FILLCELL_X1 PHY_794 ();
 FILLCELL_X1 PHY_795 ();
 FILLCELL_X1 PHY_796 ();
 FILLCELL_X1 PHY_797 ();
 FILLCELL_X1 PHY_798 ();
 FILLCELL_X1 PHY_799 ();
 FILLCELL_X1 PHY_8 ();
 FILLCELL_X1 PHY_80 ();
 FILLCELL_X1 PHY_800 ();
 FILLCELL_X1 PHY_801 ();
 FILLCELL_X1 PHY_802 ();
 FILLCELL_X1 PHY_803 ();
 FILLCELL_X1 PHY_804 ();
 FILLCELL_X1 PHY_805 ();
 FILLCELL_X1 PHY_806 ();
 FILLCELL_X1 PHY_807 ();
 FILLCELL_X1 PHY_808 ();
 FILLCELL_X1 PHY_809 ();
 FILLCELL_X1 PHY_81 ();
 FILLCELL_X1 PHY_810 ();
 FILLCELL_X1 PHY_811 ();
 FILLCELL_X1 PHY_812 ();
 FILLCELL_X1 PHY_813 ();
 FILLCELL_X1 PHY_814 ();
 FILLCELL_X1 PHY_815 ();
 FILLCELL_X1 PHY_816 ();
 FILLCELL_X1 PHY_817 ();
 FILLCELL_X1 PHY_818 ();
 FILLCELL_X1 PHY_819 ();
 FILLCELL_X1 PHY_82 ();
 FILLCELL_X1 PHY_820 ();
 FILLCELL_X1 PHY_821 ();
 FILLCELL_X1 PHY_822 ();
 FILLCELL_X1 PHY_823 ();
 FILLCELL_X1 PHY_824 ();
 FILLCELL_X1 PHY_825 ();
 FILLCELL_X1 PHY_826 ();
 FILLCELL_X1 PHY_827 ();
 FILLCELL_X1 PHY_828 ();
 FILLCELL_X1 PHY_829 ();
 FILLCELL_X1 PHY_83 ();
 FILLCELL_X1 PHY_830 ();
 FILLCELL_X1 PHY_831 ();
 FILLCELL_X1 PHY_832 ();
 FILLCELL_X1 PHY_833 ();
 FILLCELL_X1 PHY_834 ();
 FILLCELL_X1 PHY_835 ();
 FILLCELL_X1 PHY_836 ();
 FILLCELL_X1 PHY_837 ();
 FILLCELL_X1 PHY_838 ();
 FILLCELL_X1 PHY_839 ();
 FILLCELL_X1 PHY_84 ();
 FILLCELL_X1 PHY_840 ();
 FILLCELL_X1 PHY_841 ();
 FILLCELL_X1 PHY_842 ();
 FILLCELL_X1 PHY_843 ();
 FILLCELL_X1 PHY_844 ();
 FILLCELL_X1 PHY_845 ();
 FILLCELL_X1 PHY_846 ();
 FILLCELL_X1 PHY_847 ();
 FILLCELL_X1 PHY_848 ();
 FILLCELL_X1 PHY_849 ();
 FILLCELL_X1 PHY_85 ();
 FILLCELL_X1 PHY_850 ();
 FILLCELL_X1 PHY_851 ();
 FILLCELL_X1 PHY_852 ();
 FILLCELL_X1 PHY_853 ();
 FILLCELL_X1 PHY_854 ();
 FILLCELL_X1 PHY_855 ();
 FILLCELL_X1 PHY_856 ();
 FILLCELL_X1 PHY_857 ();
 FILLCELL_X1 PHY_858 ();
 FILLCELL_X1 PHY_859 ();
 FILLCELL_X1 PHY_86 ();
 FILLCELL_X1 PHY_860 ();
 FILLCELL_X1 PHY_861 ();
 FILLCELL_X1 PHY_862 ();
 FILLCELL_X1 PHY_863 ();
 FILLCELL_X1 PHY_864 ();
 FILLCELL_X1 PHY_865 ();
 FILLCELL_X1 PHY_866 ();
 FILLCELL_X1 PHY_867 ();
 FILLCELL_X1 PHY_868 ();
 FILLCELL_X1 PHY_869 ();
 FILLCELL_X1 PHY_87 ();
 FILLCELL_X1 PHY_870 ();
 FILLCELL_X1 PHY_871 ();
 FILLCELL_X1 PHY_872 ();
 FILLCELL_X1 PHY_873 ();
 FILLCELL_X1 PHY_874 ();
 FILLCELL_X1 PHY_875 ();
 FILLCELL_X1 PHY_876 ();
 FILLCELL_X1 PHY_877 ();
 FILLCELL_X1 PHY_878 ();
 FILLCELL_X1 PHY_879 ();
 FILLCELL_X1 PHY_88 ();
 FILLCELL_X1 PHY_880 ();
 FILLCELL_X1 PHY_881 ();
 FILLCELL_X1 PHY_882 ();
 FILLCELL_X1 PHY_883 ();
 FILLCELL_X1 PHY_884 ();
 FILLCELL_X1 PHY_885 ();
 FILLCELL_X1 PHY_886 ();
 FILLCELL_X1 PHY_887 ();
 FILLCELL_X1 PHY_888 ();
 FILLCELL_X1 PHY_889 ();
 FILLCELL_X1 PHY_89 ();
 FILLCELL_X1 PHY_890 ();
 FILLCELL_X1 PHY_891 ();
 FILLCELL_X1 PHY_892 ();
 FILLCELL_X1 PHY_893 ();
 FILLCELL_X1 PHY_894 ();
 FILLCELL_X1 PHY_895 ();
 FILLCELL_X1 PHY_896 ();
 FILLCELL_X1 PHY_897 ();
 FILLCELL_X1 PHY_898 ();
 FILLCELL_X1 PHY_899 ();
 FILLCELL_X1 PHY_9 ();
 FILLCELL_X1 PHY_90 ();
 FILLCELL_X1 PHY_900 ();
 FILLCELL_X1 PHY_901 ();
 FILLCELL_X1 PHY_902 ();
 FILLCELL_X1 PHY_903 ();
 FILLCELL_X1 PHY_904 ();
 FILLCELL_X1 PHY_905 ();
 FILLCELL_X1 PHY_906 ();
 FILLCELL_X1 PHY_907 ();
 FILLCELL_X1 PHY_908 ();
 FILLCELL_X1 PHY_909 ();
 FILLCELL_X1 PHY_91 ();
 FILLCELL_X1 PHY_910 ();
 FILLCELL_X1 PHY_911 ();
 FILLCELL_X1 PHY_912 ();
 FILLCELL_X1 PHY_913 ();
 FILLCELL_X1 PHY_914 ();
 FILLCELL_X1 PHY_915 ();
 FILLCELL_X1 PHY_916 ();
 FILLCELL_X1 PHY_917 ();
 FILLCELL_X1 PHY_918 ();
 FILLCELL_X1 PHY_919 ();
 FILLCELL_X1 PHY_92 ();
 FILLCELL_X1 PHY_920 ();
 FILLCELL_X1 PHY_921 ();
 FILLCELL_X1 PHY_922 ();
 FILLCELL_X1 PHY_923 ();
 FILLCELL_X1 PHY_924 ();
 FILLCELL_X1 PHY_925 ();
 FILLCELL_X1 PHY_926 ();
 FILLCELL_X1 PHY_927 ();
 FILLCELL_X1 PHY_928 ();
 FILLCELL_X1 PHY_929 ();
 FILLCELL_X1 PHY_93 ();
 FILLCELL_X1 PHY_930 ();
 FILLCELL_X1 PHY_931 ();
 FILLCELL_X1 PHY_932 ();
 FILLCELL_X1 PHY_933 ();
 FILLCELL_X1 PHY_934 ();
 FILLCELL_X1 PHY_935 ();
 FILLCELL_X1 PHY_936 ();
 FILLCELL_X1 PHY_937 ();
 FILLCELL_X1 PHY_938 ();
 FILLCELL_X1 PHY_939 ();
 FILLCELL_X1 PHY_94 ();
 FILLCELL_X1 PHY_940 ();
 FILLCELL_X1 PHY_941 ();
 FILLCELL_X1 PHY_942 ();
 FILLCELL_X1 PHY_943 ();
 FILLCELL_X1 PHY_944 ();
 FILLCELL_X1 PHY_945 ();
 FILLCELL_X1 PHY_946 ();
 FILLCELL_X1 PHY_947 ();
 FILLCELL_X1 PHY_948 ();
 FILLCELL_X1 PHY_949 ();
 FILLCELL_X1 PHY_95 ();
 FILLCELL_X1 PHY_950 ();
 FILLCELL_X1 PHY_951 ();
 FILLCELL_X1 PHY_952 ();
 FILLCELL_X1 PHY_953 ();
 FILLCELL_X1 PHY_954 ();
 FILLCELL_X1 PHY_955 ();
 FILLCELL_X1 PHY_956 ();
 FILLCELL_X1 PHY_957 ();
 FILLCELL_X1 PHY_958 ();
 FILLCELL_X1 PHY_959 ();
 FILLCELL_X1 PHY_96 ();
 FILLCELL_X1 PHY_960 ();
 FILLCELL_X1 PHY_961 ();
 FILLCELL_X1 PHY_962 ();
 FILLCELL_X1 PHY_963 ();
 FILLCELL_X1 PHY_97 ();
 FILLCELL_X1 PHY_98 ();
 FILLCELL_X1 PHY_99 ();
 INV_X1 _17655_ (.A(_01330_),
    .ZN(_03727_));
 BUF_X2 _17656_ (.A(_03727_),
    .Z(_03738_));
 BUF_X2 _17657_ (.A(_03738_),
    .Z(_03749_));
 AND2_X1 _17658_ (.A1(_17063_),
    .A2(_17064_),
    .ZN(_03760_));
 INV_X1 _17659_ (.A(_03760_),
    .ZN(_03771_));
 INV_X1 _17660_ (.A(_17065_),
    .ZN(_03782_));
 OAI21_X1 _17661_ (.A(_03749_),
    .B1(_03771_),
    .B2(_03782_),
    .ZN(_01186_));
 AND2_X1 _17662_ (.A1(_03760_),
    .A2(_17065_),
    .ZN(_03803_));
 INV_X1 _17663_ (.A(_17066_),
    .ZN(_03814_));
 NAND2_X1 _17664_ (.A1(_03803_),
    .A2(_03814_),
    .ZN(_03825_));
 BUF_X2 _17665_ (.A(_01330_),
    .Z(_03836_));
 BUF_X2 _17666_ (.A(_03836_),
    .Z(_03847_));
 NOR2_X1 _17667_ (.A1(_01330_),
    .A2(_17063_),
    .ZN(_01194_));
 INV_X1 _17668_ (.A(_17064_),
    .ZN(_03868_));
 AND2_X1 _17669_ (.A1(_01194_),
    .A2(_03868_),
    .ZN(_03879_));
 INV_X1 _17670_ (.A(_03879_),
    .ZN(_03890_));
 OAI22_X1 _17671_ (.A1(_03825_),
    .A2(_03847_),
    .B1(_03890_),
    .B2(_17065_),
    .ZN(_01187_));
 XNOR2_X1 _17672_ (.A(_03803_),
    .B(_03814_),
    .ZN(_03911_));
 XNOR2_X1 _17673_ (.A(_03760_),
    .B(_03782_),
    .ZN(_03922_));
 BUF_X2 _17674_ (.A(_03727_),
    .Z(_03933_));
 NAND3_X1 _17675_ (.A1(_03933_),
    .A2(_03868_),
    .A3(_17063_),
    .ZN(_03944_));
 OR3_X1 _17676_ (.A1(_03911_),
    .A2(_03922_),
    .A3(_03944_),
    .ZN(_03955_));
 INV_X1 _17677_ (.A(_03922_),
    .ZN(_03966_));
 NAND3_X1 _17678_ (.A1(_03911_),
    .A2(_03966_),
    .A3(_03879_),
    .ZN(_03977_));
 NAND2_X1 _17679_ (.A1(_03955_),
    .A2(_03977_),
    .ZN(_01188_));
 OR4_X1 _17680_ (.A1(_17063_),
    .A2(_03868_),
    .A3(_17065_),
    .A4(_17066_),
    .ZN(_03997_));
 AOI21_X1 _17681_ (.A(_03847_),
    .B1(_03825_),
    .B2(_03997_),
    .ZN(_01189_));
 NAND4_X1 _17682_ (.A1(_03749_),
    .A2(_03814_),
    .A3(_17063_),
    .A4(_17064_),
    .ZN(_04018_));
 NAND2_X1 _17683_ (.A1(_03977_),
    .A2(_04018_),
    .ZN(_01190_));
 NAND2_X1 _17684_ (.A1(_03922_),
    .A2(_03814_),
    .ZN(_04039_));
 OAI21_X1 _17685_ (.A(_03977_),
    .B1(_03890_),
    .B2(_04039_),
    .ZN(_01191_));
 NOR2_X1 _17686_ (.A1(_04039_),
    .A2(_03944_),
    .ZN(_01192_));
 AND4_X1 _17687_ (.A1(_17064_),
    .A2(_03922_),
    .A3(_03814_),
    .A4(_01194_),
    .ZN(_01193_));
 NOR2_X1 _17688_ (.A1(_17063_),
    .A2(_17064_),
    .ZN(_04080_));
 NOR3_X1 _17689_ (.A1(_03760_),
    .A2(_04080_),
    .A3(_03847_),
    .ZN(_01195_));
 AOI21_X1 _17690_ (.A(_01186_),
    .B1(_03782_),
    .B2(_03771_),
    .ZN(_01196_));
 AND2_X1 _17691_ (.A1(_03911_),
    .A2(_03749_),
    .ZN(_01197_));
 BUF_X2 _17692_ (.A(_17067_),
    .Z(_04121_));
 BUF_X2 _17693_ (.A(_04121_),
    .Z(_04132_));
 XOR2_X1 _17694_ (.A(_04132_),
    .B(_16935_),
    .Z(_04143_));
 INV_X1 _17695_ (.A(_16758_),
    .ZN(_04154_));
 AND2_X1 _17696_ (.A1(_04154_),
    .A2(_16757_),
    .ZN(_04165_));
 INV_X1 _17697_ (.A(_16756_),
    .ZN(_04176_));
 NOR2_X1 _17698_ (.A1(_04176_),
    .A2(_16755_),
    .ZN(_04187_));
 AND2_X1 _17699_ (.A1(_04165_),
    .A2(_04187_),
    .ZN(_04198_));
 CLKBUF_X2 _17700_ (.A(_04198_),
    .Z(_04209_));
 INV_X1 _17701_ (.A(_16753_),
    .ZN(_04220_));
 NOR2_X2 _17702_ (.A1(_04220_),
    .A2(_16754_),
    .ZN(_04231_));
 INV_X2 _17703_ (.A(_16752_),
    .ZN(_04242_));
 NOR2_X2 _17704_ (.A1(_04242_),
    .A2(_16751_),
    .ZN(_04253_));
 AND2_X2 _17705_ (.A1(_04231_),
    .A2(_04253_),
    .ZN(_04263_));
 AND2_X1 _17706_ (.A1(_04209_),
    .A2(_04263_),
    .ZN(_04274_));
 INV_X1 _17707_ (.A(_04274_),
    .ZN(_04285_));
 AND2_X1 _17708_ (.A1(_04231_),
    .A2(_04242_),
    .ZN(_04296_));
 BUF_X2 _17709_ (.A(_04296_),
    .Z(_04307_));
 NAND2_X1 _17710_ (.A1(_04209_),
    .A2(_04307_),
    .ZN(_04318_));
 AND2_X2 _17711_ (.A1(_16752_),
    .A2(_16751_),
    .ZN(_04329_));
 AND2_X2 _17712_ (.A1(_04231_),
    .A2(_04329_),
    .ZN(_04340_));
 NAND2_X1 _17713_ (.A1(_04209_),
    .A2(_04340_),
    .ZN(_04351_));
 AND3_X1 _17714_ (.A1(_04285_),
    .A2(_04318_),
    .A3(_04351_),
    .ZN(_04362_));
 AND2_X1 _17715_ (.A1(_16753_),
    .A2(_16754_),
    .ZN(_04373_));
 CLKBUF_X2 _17716_ (.A(_04373_),
    .Z(_04384_));
 AND2_X2 _17717_ (.A1(_04253_),
    .A2(_04384_),
    .ZN(_04395_));
 AND2_X1 _17718_ (.A1(_04198_),
    .A2(_04395_),
    .ZN(_04406_));
 INV_X1 _17719_ (.A(_04406_),
    .ZN(_04417_));
 NOR2_X1 _17720_ (.A1(_16753_),
    .A2(_16754_),
    .ZN(_04428_));
 CLKBUF_X2 _17721_ (.A(_04428_),
    .Z(_04439_));
 AND2_X1 _17722_ (.A1(_04439_),
    .A2(_16751_),
    .ZN(_04450_));
 CLKBUF_X2 _17723_ (.A(_04165_),
    .Z(_04461_));
 CLKBUF_X2 _17724_ (.A(_04187_),
    .Z(_04472_));
 NAND3_X1 _17725_ (.A1(_04450_),
    .A2(_04461_),
    .A3(_04472_),
    .ZN(_04483_));
 BUF_X2 _17726_ (.A(_04209_),
    .Z(_04494_));
 INV_X1 _17727_ (.A(_16754_),
    .ZN(_04504_));
 NOR2_X1 _17728_ (.A1(_04504_),
    .A2(_16753_),
    .ZN(_04515_));
 NAND2_X2 _17729_ (.A1(_04515_),
    .A2(_04242_),
    .ZN(_04526_));
 INV_X2 _17730_ (.A(_04526_),
    .ZN(_04537_));
 AND2_X1 _17731_ (.A1(_04515_),
    .A2(_04329_),
    .ZN(_04548_));
 CLKBUF_X2 _17732_ (.A(_04548_),
    .Z(_04559_));
 OAI21_X1 _17733_ (.A(_04494_),
    .B1(_04537_),
    .B2(_04559_),
    .ZN(_04570_));
 NAND4_X1 _17734_ (.A1(_04362_),
    .A2(_04417_),
    .A3(_04483_),
    .A4(_04570_),
    .ZN(_04581_));
 NOR2_X2 _17735_ (.A1(_16756_),
    .A2(_16755_),
    .ZN(_04592_));
 AND2_X1 _17736_ (.A1(_04461_),
    .A2(_04592_),
    .ZN(_04603_));
 BUF_X2 _17737_ (.A(_04603_),
    .Z(_04614_));
 AND2_X1 _17738_ (.A1(_04384_),
    .A2(_04242_),
    .ZN(_04625_));
 BUF_X2 _17739_ (.A(_04625_),
    .Z(_04636_));
 OAI21_X1 _17740_ (.A(_04614_),
    .B1(_04395_),
    .B2(_04636_),
    .ZN(_04647_));
 CLKBUF_X2 _17741_ (.A(_04515_),
    .Z(_04658_));
 CLKBUF_X2 _17742_ (.A(_04658_),
    .Z(_04669_));
 CLKBUF_X2 _17743_ (.A(_16751_),
    .Z(_04680_));
 NAND4_X1 _17744_ (.A1(_04461_),
    .A2(_04669_),
    .A3(_04680_),
    .A4(_04592_),
    .ZN(_04691_));
 AND2_X1 _17745_ (.A1(_04647_),
    .A2(_04691_),
    .ZN(_04702_));
 CLKBUF_X2 _17746_ (.A(_04231_),
    .Z(_04713_));
 NOR2_X1 _17747_ (.A1(_16752_),
    .A2(_16751_),
    .ZN(_04724_));
 CLKBUF_X2 _17748_ (.A(_04724_),
    .Z(_04735_));
 AND2_X2 _17749_ (.A1(_04713_),
    .A2(_04735_),
    .ZN(_04746_));
 NAND2_X1 _17750_ (.A1(_04614_),
    .A2(_04746_),
    .ZN(_04756_));
 AND2_X1 _17751_ (.A1(_04428_),
    .A2(_04242_),
    .ZN(_04767_));
 BUF_X2 _17752_ (.A(_04767_),
    .Z(_04778_));
 INV_X1 _17753_ (.A(_04778_),
    .ZN(_04789_));
 INV_X2 _17754_ (.A(_04603_),
    .ZN(_04800_));
 OAI211_X1 _17755_ (.A(_04702_),
    .B(_04756_),
    .C1(_04789_),
    .C2(_04800_),
    .ZN(_04811_));
 AND2_X1 _17756_ (.A1(_16756_),
    .A2(_16755_),
    .ZN(_04822_));
 CLKBUF_X2 _17757_ (.A(_04822_),
    .Z(_04833_));
 AND2_X1 _17758_ (.A1(_04165_),
    .A2(_04833_),
    .ZN(_04844_));
 AND2_X1 _17759_ (.A1(_04713_),
    .A2(_16751_),
    .ZN(_04855_));
 AND2_X1 _17760_ (.A1(_04844_),
    .A2(_04855_),
    .ZN(_04866_));
 INV_X1 _17761_ (.A(_04866_),
    .ZN(_04877_));
 BUF_X2 _17762_ (.A(_04844_),
    .Z(_04888_));
 INV_X2 _17763_ (.A(_04329_),
    .ZN(_04899_));
 INV_X1 _17764_ (.A(_04373_),
    .ZN(_04910_));
 NOR2_X2 _17765_ (.A1(_04910_),
    .A2(_04735_),
    .ZN(_04921_));
 NAND3_X1 _17766_ (.A1(_04888_),
    .A2(_04899_),
    .A3(_04921_),
    .ZN(_04931_));
 NAND3_X1 _17767_ (.A1(_04559_),
    .A2(_04461_),
    .A3(_04833_),
    .ZN(_04940_));
 CLKBUF_X2 _17768_ (.A(_04439_),
    .Z(_04950_));
 BUF_X2 _17769_ (.A(_04242_),
    .Z(_04959_));
 OAI211_X1 _17770_ (.A(_04888_),
    .B(_04950_),
    .C1(_04959_),
    .C2(_04680_),
    .ZN(_04969_));
 NAND4_X1 _17771_ (.A1(_04877_),
    .A2(_04931_),
    .A3(_04940_),
    .A4(_04969_),
    .ZN(_04978_));
 AND2_X1 _17772_ (.A1(_04176_),
    .A2(_16755_),
    .ZN(_04988_));
 AND2_X1 _17773_ (.A1(_04165_),
    .A2(_04988_),
    .ZN(_04997_));
 AND2_X1 _17774_ (.A1(_04329_),
    .A2(_04439_),
    .ZN(_05007_));
 CLKBUF_X2 _17775_ (.A(_05007_),
    .Z(_05017_));
 AND2_X1 _17776_ (.A1(_04997_),
    .A2(_05017_),
    .ZN(_05026_));
 INV_X1 _17777_ (.A(_05026_),
    .ZN(_05036_));
 CLKBUF_X2 _17778_ (.A(_04997_),
    .Z(_05045_));
 AND2_X1 _17779_ (.A1(_04231_),
    .A2(_16752_),
    .ZN(_05055_));
 BUF_X2 _17780_ (.A(_05055_),
    .Z(_05064_));
 NAND2_X1 _17781_ (.A1(_05045_),
    .A2(_05064_),
    .ZN(_05073_));
 AND2_X1 _17782_ (.A1(_04658_),
    .A2(_04680_),
    .ZN(_05082_));
 AND2_X1 _17783_ (.A1(_04329_),
    .A2(_04384_),
    .ZN(_05092_));
 BUF_X2 _17784_ (.A(_05092_),
    .Z(_05096_));
 OAI21_X1 _17785_ (.A(_05045_),
    .B1(_05082_),
    .B2(_05096_),
    .ZN(_05101_));
 NAND2_X1 _17786_ (.A1(_05045_),
    .A2(_04778_),
    .ZN(_05103_));
 NAND4_X1 _17787_ (.A1(_05036_),
    .A2(_05073_),
    .A3(_05101_),
    .A4(_05103_),
    .ZN(_05106_));
 NOR4_X1 _17788_ (.A1(_04581_),
    .A2(_04811_),
    .A3(_04978_),
    .A4(_05106_),
    .ZN(_05108_));
 NOR2_X2 _17789_ (.A1(_04154_),
    .A2(_16757_),
    .ZN(_05110_));
 AND2_X1 _17790_ (.A1(_04988_),
    .A2(_05110_),
    .ZN(_05112_));
 INV_X1 _17791_ (.A(_05112_),
    .ZN(_05114_));
 INV_X1 _17792_ (.A(_16751_),
    .ZN(_05116_));
 NOR2_X1 _17793_ (.A1(_05116_),
    .A2(_16752_),
    .ZN(_05118_));
 AND2_X2 _17794_ (.A1(_05118_),
    .A2(_04439_),
    .ZN(_05120_));
 INV_X1 _17795_ (.A(_05120_),
    .ZN(_05126_));
 CLKBUF_X2 _17796_ (.A(_16752_),
    .Z(_05137_));
 AND2_X1 _17797_ (.A1(_04384_),
    .A2(_05137_),
    .ZN(_05148_));
 BUF_X2 _17798_ (.A(_05148_),
    .Z(_05159_));
 INV_X1 _17799_ (.A(_05159_),
    .ZN(_05170_));
 AOI21_X1 _17800_ (.A(_05114_),
    .B1(_05126_),
    .B2(_05170_),
    .ZN(_05181_));
 CLKBUF_X2 _17801_ (.A(_05116_),
    .Z(_05192_));
 BUF_X2 _17802_ (.A(_05192_),
    .Z(_05203_));
 CLKBUF_X2 _17803_ (.A(_05112_),
    .Z(_05214_));
 AND2_X2 _17804_ (.A1(_04428_),
    .A2(_05137_),
    .ZN(_05225_));
 AND2_X1 _17805_ (.A1(_05214_),
    .A2(_05225_),
    .ZN(_05236_));
 AOI21_X1 _17806_ (.A(_05181_),
    .B1(_05203_),
    .B2(_05236_),
    .ZN(_05247_));
 AND2_X1 _17807_ (.A1(_04472_),
    .A2(_05110_),
    .ZN(_05258_));
 AND2_X1 _17808_ (.A1(_05258_),
    .A2(_04746_),
    .ZN(_05269_));
 INV_X1 _17809_ (.A(_05269_),
    .ZN(_05280_));
 CLKBUF_X2 _17810_ (.A(_05258_),
    .Z(_05291_));
 OAI21_X1 _17811_ (.A(_05291_),
    .B1(_05096_),
    .B2(_04636_),
    .ZN(_05302_));
 CLKBUF_X2 _17812_ (.A(_05118_),
    .Z(_05313_));
 CLKBUF_X2 _17813_ (.A(_05110_),
    .Z(_05324_));
 NAND4_X1 _17814_ (.A1(_05313_),
    .A2(_04669_),
    .A3(_04472_),
    .A4(_05324_),
    .ZN(_05335_));
 NAND3_X1 _17815_ (.A1(_05280_),
    .A2(_05302_),
    .A3(_05335_),
    .ZN(_05346_));
 INV_X1 _17816_ (.A(_04231_),
    .ZN(_05357_));
 CLKBUF_X2 _17817_ (.A(_04253_),
    .Z(_05368_));
 NOR2_X1 _17818_ (.A1(_05357_),
    .A2(_05368_),
    .ZN(_05379_));
 AND2_X1 _17819_ (.A1(_05110_),
    .A2(_04822_),
    .ZN(_05390_));
 BUF_X2 _17820_ (.A(_05390_),
    .Z(_05401_));
 AND2_X1 _17821_ (.A1(_05379_),
    .A2(_05401_),
    .ZN(_05412_));
 INV_X1 _17822_ (.A(_05390_),
    .ZN(_05423_));
 INV_X1 _17823_ (.A(_05225_),
    .ZN(_05434_));
 AND2_X1 _17824_ (.A1(_04428_),
    .A2(_04735_),
    .ZN(_05445_));
 INV_X1 _17825_ (.A(_05445_),
    .ZN(_05456_));
 AOI21_X1 _17826_ (.A(_05423_),
    .B1(_05434_),
    .B2(_05456_),
    .ZN(_05467_));
 AND2_X1 _17827_ (.A1(_04384_),
    .A2(_04735_),
    .ZN(_05478_));
 AND3_X1 _17828_ (.A1(_05478_),
    .A2(_04833_),
    .A3(_05324_),
    .ZN(_05489_));
 NOR4_X1 _17829_ (.A1(_05346_),
    .A2(_05412_),
    .A3(_05467_),
    .A4(_05489_),
    .ZN(_05500_));
 AND2_X2 _17830_ (.A1(_05110_),
    .A2(_04592_),
    .ZN(_05511_));
 BUF_X2 _17831_ (.A(_05511_),
    .Z(_05522_));
 AND2_X1 _17832_ (.A1(_04439_),
    .A2(_05116_),
    .ZN(_05533_));
 OAI21_X1 _17833_ (.A(_05522_),
    .B1(_05379_),
    .B2(_05533_),
    .ZN(_05544_));
 OAI21_X1 _17834_ (.A(_05522_),
    .B1(_04921_),
    .B2(_05082_),
    .ZN(_05555_));
 AND4_X1 _17835_ (.A1(_05247_),
    .A2(_05500_),
    .A3(_05544_),
    .A4(_05555_),
    .ZN(_05566_));
 AND2_X1 _17836_ (.A1(_16758_),
    .A2(_16757_),
    .ZN(_05577_));
 AND2_X1 _17837_ (.A1(_04988_),
    .A2(_05577_),
    .ZN(_05588_));
 AND2_X2 _17838_ (.A1(_04253_),
    .A2(_04515_),
    .ZN(_05599_));
 AND2_X1 _17839_ (.A1(_05588_),
    .A2(_05599_),
    .ZN(_05610_));
 INV_X1 _17840_ (.A(_05610_),
    .ZN(_05621_));
 CLKBUF_X2 _17841_ (.A(_05588_),
    .Z(_05632_));
 NAND2_X1 _17842_ (.A1(_05632_),
    .A2(_04559_),
    .ZN(_05643_));
 INV_X1 _17843_ (.A(_05632_),
    .ZN(_05654_));
 OAI211_X1 _17844_ (.A(_05621_),
    .B(_05643_),
    .C1(_05654_),
    .C2(_04526_),
    .ZN(_05665_));
 AND2_X2 _17845_ (.A1(_04253_),
    .A2(_04439_),
    .ZN(_05676_));
 CLKBUF_X2 _17846_ (.A(_04988_),
    .Z(_05687_));
 AND3_X1 _17847_ (.A1(_05676_),
    .A2(_05687_),
    .A3(_05577_),
    .ZN(_05698_));
 AND2_X1 _17848_ (.A1(_04231_),
    .A2(_05118_),
    .ZN(_05709_));
 AND3_X1 _17849_ (.A1(_05709_),
    .A2(_05687_),
    .A3(_05577_),
    .ZN(_05720_));
 OR2_X1 _17850_ (.A1(_05698_),
    .A2(_05720_),
    .ZN(_05731_));
 AND3_X1 _17851_ (.A1(_05632_),
    .A2(_04899_),
    .A3(_04921_),
    .ZN(_05742_));
 NOR3_X1 _17852_ (.A1(_05665_),
    .A2(_05731_),
    .A3(_05742_),
    .ZN(_05753_));
 AND2_X1 _17853_ (.A1(_05577_),
    .A2(_04592_),
    .ZN(_05764_));
 BUF_X2 _17854_ (.A(_05764_),
    .Z(_05775_));
 BUF_X2 _17855_ (.A(_05775_),
    .Z(_05786_));
 CLKBUF_X2 _17856_ (.A(_04384_),
    .Z(_05797_));
 AND3_X1 _17857_ (.A1(_05786_),
    .A2(_05368_),
    .A3(_05797_),
    .ZN(_05808_));
 AND2_X1 _17858_ (.A1(_05082_),
    .A2(_05786_),
    .ZN(_05819_));
 AND3_X1 _17859_ (.A1(_05775_),
    .A2(_05192_),
    .A3(_05225_),
    .ZN(_05830_));
 AND2_X1 _17860_ (.A1(_04636_),
    .A2(_05775_),
    .ZN(_05841_));
 NOR4_X1 _17861_ (.A1(_05808_),
    .A2(_05819_),
    .A3(_05830_),
    .A4(_05841_),
    .ZN(_05852_));
 BUF_X2 _17862_ (.A(_04658_),
    .Z(_05863_));
 BUF_X2 _17863_ (.A(_05577_),
    .Z(_05874_));
 NAND4_X1 _17864_ (.A1(_05863_),
    .A2(_04472_),
    .A3(_04735_),
    .A4(_05874_),
    .ZN(_05885_));
 AND2_X1 _17865_ (.A1(_04472_),
    .A2(_05577_),
    .ZN(_05896_));
 BUF_X2 _17866_ (.A(_05896_),
    .Z(_05907_));
 INV_X1 _17867_ (.A(_05007_),
    .ZN(_05918_));
 NAND2_X1 _17868_ (.A1(_05918_),
    .A2(_05456_),
    .ZN(_05929_));
 OAI21_X1 _17869_ (.A(_05907_),
    .B1(_05929_),
    .B2(_04307_),
    .ZN(_05940_));
 OAI211_X1 _17870_ (.A(_05907_),
    .B(_04669_),
    .C1(_05368_),
    .C2(_04329_),
    .ZN(_05951_));
 AND2_X1 _17871_ (.A1(_04384_),
    .A2(_16751_),
    .ZN(_05962_));
 AND2_X1 _17872_ (.A1(_05896_),
    .A2(_05962_),
    .ZN(_05973_));
 INV_X1 _17873_ (.A(_05973_),
    .ZN(_05984_));
 AND4_X1 _17874_ (.A1(_05885_),
    .A2(_05940_),
    .A3(_05951_),
    .A4(_05984_),
    .ZN(_05995_));
 AND2_X1 _17875_ (.A1(_04822_),
    .A2(_05577_),
    .ZN(_06006_));
 CLKBUF_X2 _17876_ (.A(_06006_),
    .Z(_06017_));
 AND2_X1 _17877_ (.A1(_04746_),
    .A2(_06017_),
    .ZN(_06028_));
 INV_X1 _17878_ (.A(_06028_),
    .ZN(_06039_));
 NAND2_X1 _17879_ (.A1(_06017_),
    .A2(_05225_),
    .ZN(_06050_));
 NAND2_X1 _17880_ (.A1(_05120_),
    .A2(_06017_),
    .ZN(_06061_));
 OAI211_X1 _17881_ (.A(_06017_),
    .B(_16754_),
    .C1(_04220_),
    .C2(_05368_),
    .ZN(_06072_));
 AND4_X1 _17882_ (.A1(_06039_),
    .A2(_06050_),
    .A3(_06061_),
    .A4(_06072_),
    .ZN(_06083_));
 AND4_X1 _17883_ (.A1(_05753_),
    .A2(_05852_),
    .A3(_05995_),
    .A4(_06083_),
    .ZN(_06094_));
 INV_X1 _17884_ (.A(_04548_),
    .ZN(_06105_));
 AND2_X1 _17885_ (.A1(_04658_),
    .A2(_04735_),
    .ZN(_06116_));
 INV_X1 _17886_ (.A(_06116_),
    .ZN(_06127_));
 NAND2_X1 _17887_ (.A1(_06105_),
    .A2(_06127_),
    .ZN(_06138_));
 NOR2_X2 _17888_ (.A1(_16758_),
    .A2(_16757_),
    .ZN(_06149_));
 AND2_X2 _17889_ (.A1(_05687_),
    .A2(_06149_),
    .ZN(_06160_));
 CLKBUF_X2 _17890_ (.A(_06160_),
    .Z(_06171_));
 AND2_X1 _17891_ (.A1(_06138_),
    .A2(_06171_),
    .ZN(_06182_));
 INV_X1 _17892_ (.A(_06182_),
    .ZN(_06193_));
 NAND3_X1 _17893_ (.A1(_05225_),
    .A2(_06149_),
    .A3(_05687_),
    .ZN(_06204_));
 INV_X1 _17894_ (.A(_06160_),
    .ZN(_06215_));
 AND2_X1 _17895_ (.A1(_04899_),
    .A2(_04231_),
    .ZN(_06226_));
 INV_X1 _17896_ (.A(_04724_),
    .ZN(_06236_));
 AND2_X1 _17897_ (.A1(_06226_),
    .A2(_06236_),
    .ZN(_06238_));
 INV_X1 _17898_ (.A(_06238_),
    .ZN(_06248_));
 OAI211_X1 _17899_ (.A(_06193_),
    .B(_06204_),
    .C1(_06215_),
    .C2(_06248_),
    .ZN(_06259_));
 AND2_X2 _17900_ (.A1(_06149_),
    .A2(_04592_),
    .ZN(_06270_));
 CLKBUF_X2 _17901_ (.A(_06270_),
    .Z(_06281_));
 NAND3_X1 _17902_ (.A1(_04921_),
    .A2(_04899_),
    .A3(_06281_),
    .ZN(_06292_));
 BUF_X2 _17903_ (.A(_04713_),
    .Z(_06303_));
 BUF_X2 _17904_ (.A(_05137_),
    .Z(_06314_));
 CLKBUF_X2 _17905_ (.A(_04680_),
    .Z(_06325_));
 OAI211_X1 _17906_ (.A(_06281_),
    .B(_06303_),
    .C1(_06314_),
    .C2(_06325_),
    .ZN(_06336_));
 OAI211_X1 _17907_ (.A(_06281_),
    .B(_05863_),
    .C1(_06314_),
    .C2(_04680_),
    .ZN(_06347_));
 NAND2_X1 _17908_ (.A1(_06281_),
    .A2(_05225_),
    .ZN(_06358_));
 NAND4_X1 _17909_ (.A1(_06292_),
    .A2(_06336_),
    .A3(_06347_),
    .A4(_06358_),
    .ZN(_06369_));
 AND2_X1 _17910_ (.A1(_04472_),
    .A2(_06149_),
    .ZN(_06380_));
 BUF_X2 _17911_ (.A(_06380_),
    .Z(_06391_));
 INV_X1 _17912_ (.A(_04439_),
    .ZN(_06402_));
 NOR2_X1 _17913_ (.A1(_06402_),
    .A2(_04329_),
    .ZN(_06413_));
 AND2_X1 _17914_ (.A1(_06391_),
    .A2(_06413_),
    .ZN(_06424_));
 INV_X1 _17915_ (.A(_06424_),
    .ZN(_06435_));
 BUF_X2 _17916_ (.A(_06391_),
    .Z(_06446_));
 NAND4_X1 _17917_ (.A1(_06446_),
    .A2(_06303_),
    .A3(_04899_),
    .A4(_06236_),
    .ZN(_06457_));
 AND2_X1 _17918_ (.A1(_06236_),
    .A2(_04515_),
    .ZN(_06468_));
 NAND2_X1 _17919_ (.A1(_06468_),
    .A2(_06446_),
    .ZN(_06479_));
 BUF_X2 _17920_ (.A(_05478_),
    .Z(_06490_));
 OAI21_X1 _17921_ (.A(_06446_),
    .B1(_06490_),
    .B2(_05159_),
    .ZN(_06501_));
 NAND4_X1 _17922_ (.A1(_06435_),
    .A2(_06457_),
    .A3(_06479_),
    .A4(_06501_),
    .ZN(_06512_));
 NAND2_X1 _17923_ (.A1(_06236_),
    .A2(_04439_),
    .ZN(_06523_));
 INV_X1 _17924_ (.A(_06523_),
    .ZN(_06534_));
 AND2_X1 _17925_ (.A1(_04822_),
    .A2(_06149_),
    .ZN(_06545_));
 CLKBUF_X2 _17926_ (.A(_06545_),
    .Z(_06556_));
 BUF_X2 _17927_ (.A(_06556_),
    .Z(_06567_));
 NAND2_X1 _17928_ (.A1(_06534_),
    .A2(_06567_),
    .ZN(_06578_));
 OAI211_X1 _17929_ (.A(_06567_),
    .B(_05797_),
    .C1(_04959_),
    .C2(_04680_),
    .ZN(_06589_));
 NAND2_X1 _17930_ (.A1(_06116_),
    .A2(_06567_),
    .ZN(_06600_));
 NAND3_X1 _17931_ (.A1(_06567_),
    .A2(_06303_),
    .A3(_05368_),
    .ZN(_06611_));
 NAND4_X1 _17932_ (.A1(_06578_),
    .A2(_06589_),
    .A3(_06600_),
    .A4(_06611_),
    .ZN(_06622_));
 NOR4_X1 _17933_ (.A1(_06259_),
    .A2(_06369_),
    .A3(_06512_),
    .A4(_06622_),
    .ZN(_06633_));
 NAND4_X1 _17934_ (.A1(_05108_),
    .A2(_05566_),
    .A3(_06094_),
    .A4(_06633_),
    .ZN(_06644_));
 OAI21_X1 _17935_ (.A(_04504_),
    .B1(_06236_),
    .B2(_16753_),
    .ZN(_06655_));
 AND3_X1 _17936_ (.A1(_06149_),
    .A2(_04592_),
    .A3(_04504_),
    .ZN(_06666_));
 AND2_X1 _17937_ (.A1(_06655_),
    .A2(_06666_),
    .ZN(_06672_));
 NOR2_X2 _17938_ (.A1(_06644_),
    .A2(_06672_),
    .ZN(_06677_));
 NOR2_X1 _17939_ (.A1(_16716_),
    .A2(_16715_),
    .ZN(_06688_));
 CLKBUF_X2 _17940_ (.A(_06688_),
    .Z(_06699_));
 NOR2_X1 _17941_ (.A1(_16718_),
    .A2(_16717_),
    .ZN(_06710_));
 AND2_X1 _17942_ (.A1(_06699_),
    .A2(_06710_),
    .ZN(_06721_));
 BUF_X2 _17943_ (.A(_06721_),
    .Z(_06732_));
 NOR2_X2 _17944_ (.A1(_16713_),
    .A2(_16714_),
    .ZN(_06743_));
 CLKBUF_X2 _17945_ (.A(_16712_),
    .Z(_06754_));
 AND2_X1 _17946_ (.A1(_06743_),
    .A2(_06754_),
    .ZN(_06765_));
 BUF_X2 _17947_ (.A(_06765_),
    .Z(_06776_));
 AND2_X1 _17948_ (.A1(_06732_),
    .A2(_06776_),
    .ZN(_06787_));
 INV_X1 _17949_ (.A(_16717_),
    .ZN(_06798_));
 AND2_X1 _17950_ (.A1(_06798_),
    .A2(_16718_),
    .ZN(_06809_));
 AND2_X1 _17951_ (.A1(_16716_),
    .A2(_16715_),
    .ZN(_06820_));
 AND2_X1 _17952_ (.A1(_06809_),
    .A2(_06820_),
    .ZN(_06831_));
 INV_X2 _17953_ (.A(_06743_),
    .ZN(_06842_));
 INV_X1 _17954_ (.A(_16711_),
    .ZN(_06853_));
 NOR2_X1 _17955_ (.A1(_06853_),
    .A2(_16712_),
    .ZN(_06864_));
 BUF_X2 _17956_ (.A(_06864_),
    .Z(_06875_));
 NOR2_X1 _17957_ (.A1(_06842_),
    .A2(_06875_),
    .ZN(_06886_));
 AND2_X1 _17958_ (.A1(_06831_),
    .A2(_06886_),
    .ZN(_06897_));
 INV_X1 _17959_ (.A(_16713_),
    .ZN(_06908_));
 NOR2_X2 _17960_ (.A1(_06908_),
    .A2(_16714_),
    .ZN(_06919_));
 INV_X2 _17961_ (.A(_16712_),
    .ZN(_06930_));
 AND2_X1 _17962_ (.A1(_06919_),
    .A2(_06930_),
    .ZN(_06941_));
 BUF_X2 _17963_ (.A(_06941_),
    .Z(_06952_));
 INV_X1 _17964_ (.A(_16716_),
    .ZN(_06963_));
 NOR2_X2 _17965_ (.A1(_06963_),
    .A2(_16715_),
    .ZN(_06974_));
 AND2_X1 _17966_ (.A1(_16718_),
    .A2(_16717_),
    .ZN(_06985_));
 AND2_X1 _17967_ (.A1(_06974_),
    .A2(_06985_),
    .ZN(_06996_));
 CLKBUF_X2 _17968_ (.A(_06996_),
    .Z(_07007_));
 AND2_X1 _17969_ (.A1(_06952_),
    .A2(_07007_),
    .ZN(_07018_));
 NOR2_X1 _17970_ (.A1(_16712_),
    .A2(_16711_),
    .ZN(_07021_));
 AND2_X2 _17971_ (.A1(_06743_),
    .A2(_07021_),
    .ZN(_07029_));
 AND2_X1 _17972_ (.A1(_07029_),
    .A2(_06721_),
    .ZN(_07040_));
 OR4_X1 _17973_ (.A1(_06787_),
    .A2(_06897_),
    .A3(_07018_),
    .A4(_07040_),
    .ZN(_07051_));
 NOR2_X2 _17974_ (.A1(_06798_),
    .A2(_16718_),
    .ZN(_07062_));
 AND2_X1 _17975_ (.A1(_06974_),
    .A2(_07062_),
    .ZN(_07073_));
 BUF_X2 _17976_ (.A(_07073_),
    .Z(_07084_));
 BUF_X2 _17977_ (.A(_07084_),
    .Z(_07095_));
 INV_X1 _17978_ (.A(_16714_),
    .ZN(_07106_));
 NOR2_X2 _17979_ (.A1(_07106_),
    .A2(_16713_),
    .ZN(_07117_));
 INV_X1 _17980_ (.A(_07117_),
    .ZN(_07128_));
 NOR2_X2 _17981_ (.A1(_06930_),
    .A2(_16711_),
    .ZN(_07139_));
 BUF_X2 _17982_ (.A(_07139_),
    .Z(_07150_));
 CLKBUF_X2 _17983_ (.A(_06853_),
    .Z(_07161_));
 OAI22_X1 _17984_ (.A1(_07128_),
    .A2(_07150_),
    .B1(_07161_),
    .B2(_06842_),
    .ZN(_07172_));
 BUF_X1 _17985_ (.A(_06919_),
    .Z(_07183_));
 CLKBUF_X2 _17986_ (.A(_07183_),
    .Z(_07194_));
 OAI21_X1 _17987_ (.A(_07095_),
    .B1(_07172_),
    .B2(_07194_),
    .ZN(_07205_));
 AND2_X2 _17988_ (.A1(_06875_),
    .A2(_07117_),
    .ZN(_07216_));
 AND2_X1 _17989_ (.A1(_06985_),
    .A2(_06688_),
    .ZN(_07227_));
 CLKBUF_X2 _17990_ (.A(_07227_),
    .Z(_07238_));
 BUF_X2 _17991_ (.A(_07238_),
    .Z(_07249_));
 NAND2_X1 _17992_ (.A1(_07216_),
    .A2(_07249_),
    .ZN(_07260_));
 NOR2_X1 _17993_ (.A1(_07128_),
    .A2(_06875_),
    .ZN(_07271_));
 INV_X1 _17994_ (.A(_07271_),
    .ZN(_07282_));
 INV_X1 _17995_ (.A(_06996_),
    .ZN(_07293_));
 OAI211_X1 _17996_ (.A(_07205_),
    .B(_07260_),
    .C1(_07282_),
    .C2(_07293_),
    .ZN(_07304_));
 BUF_X2 _17997_ (.A(_06831_),
    .Z(_07315_));
 AND2_X1 _17998_ (.A1(_16713_),
    .A2(_16714_),
    .ZN(_07326_));
 AND2_X1 _17999_ (.A1(_07326_),
    .A2(_07021_),
    .ZN(_07337_));
 BUF_X2 _18000_ (.A(_07337_),
    .Z(_07348_));
 CLKBUF_X2 _18001_ (.A(_07326_),
    .Z(_07356_));
 AND2_X1 _18002_ (.A1(_07356_),
    .A2(_06930_),
    .ZN(_07367_));
 BUF_X2 _18003_ (.A(_07367_),
    .Z(_07378_));
 AND2_X1 _18004_ (.A1(_06820_),
    .A2(_06710_),
    .ZN(_07389_));
 BUF_X2 _18005_ (.A(_07389_),
    .Z(_07400_));
 BUF_X2 _18006_ (.A(_07400_),
    .Z(_07411_));
 AOI22_X1 _18007_ (.A1(_07315_),
    .A2(_07348_),
    .B1(_07378_),
    .B2(_07411_),
    .ZN(_07422_));
 INV_X1 _18008_ (.A(_06919_),
    .ZN(_07433_));
 NOR2_X1 _18009_ (.A1(_07433_),
    .A2(_07139_),
    .ZN(_07444_));
 AND2_X1 _18010_ (.A1(_06809_),
    .A2(_06699_),
    .ZN(_07455_));
 BUF_X2 _18011_ (.A(_07455_),
    .Z(_07466_));
 NAND2_X1 _18012_ (.A1(_07444_),
    .A2(_07466_),
    .ZN(_07477_));
 INV_X1 _18013_ (.A(_06721_),
    .ZN(_07488_));
 AND2_X1 _18014_ (.A1(_06919_),
    .A2(_06754_),
    .ZN(_07499_));
 INV_X1 _18015_ (.A(_07499_),
    .ZN(_07510_));
 OAI211_X1 _18016_ (.A(_07422_),
    .B(_07477_),
    .C1(_07488_),
    .C2(_07510_),
    .ZN(_07521_));
 AND2_X2 _18017_ (.A1(_06875_),
    .A2(_06743_),
    .ZN(_07532_));
 CLKBUF_X2 _18018_ (.A(_06985_),
    .Z(_07543_));
 CLKBUF_X2 _18019_ (.A(_06820_),
    .Z(_07554_));
 AND2_X1 _18020_ (.A1(_07543_),
    .A2(_07554_),
    .ZN(_07565_));
 BUF_X2 _18021_ (.A(_07565_),
    .Z(_07576_));
 AND2_X1 _18022_ (.A1(_16712_),
    .A2(_16711_),
    .ZN(_07587_));
 BUF_X2 _18023_ (.A(_07587_),
    .Z(_07598_));
 AND2_X2 _18024_ (.A1(_07598_),
    .A2(_07356_),
    .ZN(_07609_));
 AOI22_X1 _18025_ (.A1(_07532_),
    .A2(_07576_),
    .B1(_07609_),
    .B2(_07400_),
    .ZN(_07620_));
 AND2_X1 _18026_ (.A1(_06809_),
    .A2(_06974_),
    .ZN(_07631_));
 INV_X1 _18027_ (.A(_07631_),
    .ZN(_07641_));
 AND2_X1 _18028_ (.A1(_06919_),
    .A2(_07021_),
    .ZN(_07652_));
 INV_X1 _18029_ (.A(_07652_),
    .ZN(_07663_));
 AND2_X1 _18030_ (.A1(_07062_),
    .A2(_06820_),
    .ZN(_07674_));
 INV_X1 _18031_ (.A(_07674_),
    .ZN(_07685_));
 AND2_X1 _18032_ (.A1(_06743_),
    .A2(_06930_),
    .ZN(_07696_));
 INV_X1 _18033_ (.A(_07696_),
    .ZN(_07707_));
 OAI221_X1 _18034_ (.A(_07620_),
    .B1(_07641_),
    .B2(_07663_),
    .C1(_07685_),
    .C2(_07707_),
    .ZN(_07718_));
 NOR4_X1 _18035_ (.A1(_07051_),
    .A2(_07304_),
    .A3(_07521_),
    .A4(_07718_),
    .ZN(_07729_));
 INV_X1 _18036_ (.A(_07356_),
    .ZN(_07740_));
 NOR2_X1 _18037_ (.A1(_07740_),
    .A2(_07598_),
    .ZN(_07751_));
 AND2_X2 _18038_ (.A1(_07139_),
    .A2(_06743_),
    .ZN(_07762_));
 OAI21_X1 _18039_ (.A(_07249_),
    .B1(_07751_),
    .B2(_07762_),
    .ZN(_07773_));
 AND2_X1 _18040_ (.A1(_07139_),
    .A2(_06919_),
    .ZN(_07784_));
 BUF_X2 _18041_ (.A(_07784_),
    .Z(_07795_));
 AND2_X1 _18042_ (.A1(_07117_),
    .A2(_07021_),
    .ZN(_07806_));
 OAI21_X1 _18043_ (.A(_07411_),
    .B1(_07795_),
    .B2(_07806_),
    .ZN(_07817_));
 AND2_X1 _18044_ (.A1(_06974_),
    .A2(_06710_),
    .ZN(_07828_));
 BUF_X2 _18045_ (.A(_07828_),
    .Z(_07839_));
 INV_X1 _18046_ (.A(_07021_),
    .ZN(_07850_));
 AND2_X1 _18047_ (.A1(_07850_),
    .A2(_07117_),
    .ZN(_07861_));
 NOR2_X1 _18048_ (.A1(_06842_),
    .A2(_07598_),
    .ZN(_07872_));
 OAI21_X1 _18049_ (.A(_07839_),
    .B1(_07861_),
    .B2(_07872_),
    .ZN(_07883_));
 AND2_X2 _18050_ (.A1(_07062_),
    .A2(_06699_),
    .ZN(_07893_));
 BUF_X2 _18051_ (.A(_07696_),
    .Z(_07904_));
 OAI21_X1 _18052_ (.A(_07893_),
    .B1(_07652_),
    .B2(_07904_),
    .ZN(_07915_));
 NAND4_X1 _18053_ (.A1(_07773_),
    .A2(_07817_),
    .A3(_07883_),
    .A4(_07915_),
    .ZN(_07926_));
 AND2_X1 _18054_ (.A1(_07117_),
    .A2(_07587_),
    .ZN(_07937_));
 CLKBUF_X2 _18055_ (.A(_07937_),
    .Z(_07948_));
 INV_X1 _18056_ (.A(_07948_),
    .ZN(_07959_));
 INV_X1 _18057_ (.A(_07806_),
    .ZN(_07970_));
 NAND2_X1 _18058_ (.A1(_07959_),
    .A2(_07970_),
    .ZN(_07981_));
 AND2_X1 _18059_ (.A1(_06963_),
    .A2(_16715_),
    .ZN(_07992_));
 AND2_X1 _18060_ (.A1(_07992_),
    .A2(_06710_),
    .ZN(_08003_));
 BUF_X2 _18061_ (.A(_08003_),
    .Z(_08014_));
 BUF_X2 _18062_ (.A(_08014_),
    .Z(_08025_));
 AND2_X1 _18063_ (.A1(_07981_),
    .A2(_08025_),
    .ZN(_08036_));
 AND2_X2 _18064_ (.A1(_07139_),
    .A2(_07356_),
    .ZN(_08047_));
 OAI21_X1 _18065_ (.A(_07893_),
    .B1(_08047_),
    .B2(_07378_),
    .ZN(_08058_));
 BUF_X2 _18066_ (.A(_07117_),
    .Z(_08069_));
 CLKBUF_X2 _18067_ (.A(_07062_),
    .Z(_08080_));
 CLKBUF_X2 _18068_ (.A(_16711_),
    .Z(_08091_));
 CLKBUF_X2 _18069_ (.A(_08091_),
    .Z(_08102_));
 CLKBUF_X2 _18070_ (.A(_06699_),
    .Z(_08113_));
 NAND4_X1 _18071_ (.A1(_08069_),
    .A2(_08080_),
    .A3(_08102_),
    .A4(_08113_),
    .ZN(_08124_));
 NAND2_X1 _18072_ (.A1(_08058_),
    .A2(_08124_),
    .ZN(_08134_));
 AND2_X1 _18073_ (.A1(_07992_),
    .A2(_07062_),
    .ZN(_08145_));
 BUF_X2 _18074_ (.A(_08145_),
    .Z(_08156_));
 CLKBUF_X2 _18075_ (.A(_07499_),
    .Z(_08167_));
 NAND2_X1 _18076_ (.A1(_08156_),
    .A2(_08167_),
    .ZN(_08178_));
 BUF_X2 _18077_ (.A(_07992_),
    .Z(_08189_));
 BUF_X2 _18078_ (.A(_08189_),
    .Z(_08200_));
 CLKBUF_X2 _18079_ (.A(_06809_),
    .Z(_08211_));
 BUF_X2 _18080_ (.A(_08211_),
    .Z(_08222_));
 BUF_X2 _18081_ (.A(_07356_),
    .Z(_08233_));
 NAND4_X1 _18082_ (.A1(_08200_),
    .A2(_08222_),
    .A3(_06754_),
    .A4(_08233_),
    .ZN(_08244_));
 NAND4_X1 _18083_ (.A1(_08222_),
    .A2(_06754_),
    .A3(_08233_),
    .A4(_08113_),
    .ZN(_08255_));
 NAND4_X1 _18084_ (.A1(_08222_),
    .A2(_06875_),
    .A3(_08233_),
    .A4(_08113_),
    .ZN(_08266_));
 NAND4_X1 _18085_ (.A1(_08178_),
    .A2(_08244_),
    .A3(_08255_),
    .A4(_08266_),
    .ZN(_08277_));
 NOR4_X1 _18086_ (.A1(_07926_),
    .A2(_08036_),
    .A3(_08134_),
    .A4(_08277_),
    .ZN(_08288_));
 AND2_X1 _18087_ (.A1(_06919_),
    .A2(_06864_),
    .ZN(_08299_));
 BUF_X2 _18088_ (.A(_08299_),
    .Z(_08308_));
 INV_X1 _18089_ (.A(_08308_),
    .ZN(_08318_));
 INV_X1 _18090_ (.A(_07784_),
    .ZN(_08327_));
 NAND2_X1 _18091_ (.A1(_08318_),
    .A2(_08327_),
    .ZN(_08337_));
 NOR2_X1 _18092_ (.A1(_07740_),
    .A2(_06875_),
    .ZN(_08346_));
 OAI21_X1 _18093_ (.A(_07839_),
    .B1(_08337_),
    .B2(_08346_),
    .ZN(_08355_));
 AND2_X1 _18094_ (.A1(_08069_),
    .A2(_08091_),
    .ZN(_08365_));
 OR2_X1 _18095_ (.A1(_08365_),
    .A2(_07609_),
    .ZN(_08375_));
 NOR2_X2 _18096_ (.A1(_06842_),
    .A2(_07150_),
    .ZN(_08384_));
 OAI21_X1 _18097_ (.A(_08156_),
    .B1(_08375_),
    .B2(_08384_),
    .ZN(_08394_));
 BUF_X2 _18098_ (.A(_07021_),
    .Z(_08403_));
 NOR2_X1 _18099_ (.A1(_07740_),
    .A2(_08403_),
    .ZN(_08413_));
 BUF_X2 _18100_ (.A(_07674_),
    .Z(_08422_));
 INV_X1 _18101_ (.A(_07598_),
    .ZN(_08431_));
 NAND3_X1 _18102_ (.A1(_08413_),
    .A2(_08422_),
    .A3(_08431_),
    .ZN(_08441_));
 NAND2_X1 _18103_ (.A1(_07948_),
    .A2(_08422_),
    .ZN(_08447_));
 NAND2_X1 _18104_ (.A1(_08441_),
    .A2(_08447_),
    .ZN(_08448_));
 INV_X1 _18105_ (.A(_08448_),
    .ZN(_08449_));
 BUF_X2 _18106_ (.A(_07007_),
    .Z(_08450_));
 AND2_X2 _18107_ (.A1(_07587_),
    .A2(_06743_),
    .ZN(_08451_));
 INV_X1 _18108_ (.A(_08451_),
    .ZN(_08452_));
 INV_X1 _18109_ (.A(_07029_),
    .ZN(_08453_));
 NAND2_X1 _18110_ (.A1(_08452_),
    .A2(_08453_),
    .ZN(_08454_));
 AND2_X1 _18111_ (.A1(_07356_),
    .A2(_08091_),
    .ZN(_08455_));
 OAI21_X1 _18112_ (.A(_08450_),
    .B1(_08454_),
    .B2(_08455_),
    .ZN(_08456_));
 AND4_X1 _18113_ (.A1(_08355_),
    .A2(_08394_),
    .A3(_08449_),
    .A4(_08456_),
    .ZN(_08457_));
 INV_X1 _18114_ (.A(_07139_),
    .ZN(_08458_));
 BUF_X2 _18115_ (.A(_06930_),
    .Z(_08459_));
 OAI22_X1 _18116_ (.A1(_08458_),
    .A2(_07740_),
    .B1(_08459_),
    .B2(_06842_),
    .ZN(_08460_));
 BUF_X2 _18117_ (.A(_08069_),
    .Z(_08461_));
 OAI21_X1 _18118_ (.A(_07576_),
    .B1(_08460_),
    .B2(_08461_),
    .ZN(_08462_));
 BUF_X2 _18119_ (.A(_06710_),
    .Z(_08463_));
 NAND3_X1 _18120_ (.A1(_06776_),
    .A2(_08200_),
    .A3(_08463_),
    .ZN(_08464_));
 OAI21_X1 _18121_ (.A(_08025_),
    .B1(_08308_),
    .B2(_07795_),
    .ZN(_08465_));
 NAND3_X1 _18122_ (.A1(_08462_),
    .A2(_08464_),
    .A3(_08465_),
    .ZN(_08466_));
 AND2_X1 _18123_ (.A1(_07751_),
    .A2(_07850_),
    .ZN(_08467_));
 INV_X1 _18124_ (.A(_08467_),
    .ZN(_08468_));
 AOI22_X1 _18125_ (.A1(_08461_),
    .A2(_07850_),
    .B1(_07194_),
    .B2(_06875_),
    .ZN(_08469_));
 AOI21_X1 _18126_ (.A(_07488_),
    .B1(_08468_),
    .B2(_08469_),
    .ZN(_08470_));
 AND2_X1 _18127_ (.A1(_07444_),
    .A2(_06831_),
    .ZN(_08471_));
 NAND2_X1 _18128_ (.A1(_07652_),
    .A2(_07576_),
    .ZN(_08472_));
 NOR2_X2 _18129_ (.A1(_06842_),
    .A2(_08403_),
    .ZN(_08473_));
 NAND2_X1 _18130_ (.A1(_08473_),
    .A2(_07411_),
    .ZN(_08474_));
 NAND2_X1 _18131_ (.A1(_08472_),
    .A2(_08474_),
    .ZN(_08475_));
 NOR4_X1 _18132_ (.A1(_08466_),
    .A2(_08470_),
    .A3(_08471_),
    .A4(_08475_),
    .ZN(_08476_));
 AND4_X1 _18133_ (.A1(_07729_),
    .A2(_08288_),
    .A3(_08457_),
    .A4(_08476_),
    .ZN(_08477_));
 CLKBUF_X2 _18134_ (.A(_06743_),
    .Z(_08478_));
 AND2_X1 _18135_ (.A1(_08478_),
    .A2(_06853_),
    .ZN(_08479_));
 OAI21_X1 _18136_ (.A(_07466_),
    .B1(_08365_),
    .B2(_08479_),
    .ZN(_08480_));
 INV_X1 _18137_ (.A(_07238_),
    .ZN(_08481_));
 INV_X1 _18138_ (.A(_08047_),
    .ZN(_08482_));
 INV_X1 _18139_ (.A(_07095_),
    .ZN(_08483_));
 OAI221_X1 _18140_ (.A(_08480_),
    .B1(_07959_),
    .B2(_08481_),
    .C1(_08482_),
    .C2(_08483_),
    .ZN(_08484_));
 BUF_X2 _18141_ (.A(_07631_),
    .Z(_08485_));
 AND2_X1 _18142_ (.A1(_08485_),
    .A2(_07609_),
    .ZN(_08486_));
 INV_X1 _18143_ (.A(_08486_),
    .ZN(_08487_));
 OAI21_X1 _18144_ (.A(_08485_),
    .B1(_07216_),
    .B2(_07378_),
    .ZN(_08488_));
 NAND2_X1 _18145_ (.A1(_08487_),
    .A2(_08488_),
    .ZN(_08489_));
 AND2_X1 _18146_ (.A1(_07992_),
    .A2(_07543_),
    .ZN(_08490_));
 BUF_X2 _18147_ (.A(_08490_),
    .Z(_08491_));
 INV_X1 _18148_ (.A(_08491_),
    .ZN(_08492_));
 AOI21_X1 _18149_ (.A(_08461_),
    .B1(_08413_),
    .B2(_08431_),
    .ZN(_08493_));
 NOR2_X1 _18150_ (.A1(_08308_),
    .A2(_07762_),
    .ZN(_08494_));
 AOI21_X1 _18151_ (.A(_08492_),
    .B1(_08493_),
    .B2(_08494_),
    .ZN(_08495_));
 NAND4_X1 _18152_ (.A1(_08473_),
    .A2(_08200_),
    .A3(_08431_),
    .A4(_08222_),
    .ZN(_08496_));
 AND2_X1 _18153_ (.A1(_06919_),
    .A2(_08091_),
    .ZN(_08497_));
 BUF_X2 _18154_ (.A(_08497_),
    .Z(_08498_));
 NAND2_X1 _18155_ (.A1(_08422_),
    .A2(_08498_),
    .ZN(_08499_));
 OAI211_X1 _18156_ (.A(_08496_),
    .B(_08499_),
    .C1(_07685_),
    .C2(_08452_),
    .ZN(_08500_));
 NOR4_X1 _18157_ (.A1(_08484_),
    .A2(_08489_),
    .A3(_08495_),
    .A4(_08500_),
    .ZN(_08501_));
 AND2_X1 _18158_ (.A1(_08477_),
    .A2(_08501_),
    .ZN(_08502_));
 XNOR2_X1 _18159_ (.A(_06677_),
    .B(_08502_),
    .ZN(_08503_));
 INV_X1 _18160_ (.A(_16706_),
    .ZN(_08504_));
 NOR2_X1 _18161_ (.A1(_08504_),
    .A2(_16705_),
    .ZN(_08505_));
 CLKBUF_X2 _18162_ (.A(_08505_),
    .Z(_08506_));
 BUF_X2 _18163_ (.A(_16704_),
    .Z(_08507_));
 AND2_X1 _18164_ (.A1(_16703_),
    .A2(_08507_),
    .ZN(_08508_));
 BUF_X2 _18165_ (.A(_08508_),
    .Z(_08509_));
 AND2_X2 _18166_ (.A1(_08506_),
    .A2(_08509_),
    .ZN(_08510_));
 AND2_X1 _18167_ (.A1(_16710_),
    .A2(_16709_),
    .ZN(_08511_));
 NOR2_X2 _18168_ (.A1(_16708_),
    .A2(_16707_),
    .ZN(_08512_));
 AND2_X2 _18169_ (.A1(_08511_),
    .A2(_08512_),
    .ZN(_08513_));
 NAND2_X1 _18170_ (.A1(_08510_),
    .A2(_08513_),
    .ZN(_08514_));
 INV_X1 _18171_ (.A(_16705_),
    .ZN(_08515_));
 NOR2_X1 _18172_ (.A1(_08515_),
    .A2(_16706_),
    .ZN(_08516_));
 CLKBUF_X2 _18173_ (.A(_08516_),
    .Z(_08517_));
 NOR2_X1 _18174_ (.A1(_16703_),
    .A2(_16704_),
    .ZN(_08518_));
 AND2_X1 _18175_ (.A1(_08517_),
    .A2(_08518_),
    .ZN(_08519_));
 INV_X1 _18176_ (.A(_08519_),
    .ZN(_08520_));
 AND2_X2 _18177_ (.A1(_16708_),
    .A2(_16707_),
    .ZN(_08521_));
 AND2_X1 _18178_ (.A1(_08521_),
    .A2(_08511_),
    .ZN(_08522_));
 BUF_X2 _18179_ (.A(_08522_),
    .Z(_08523_));
 INV_X1 _18180_ (.A(_08523_),
    .ZN(_08524_));
 INV_X1 _18181_ (.A(_16703_),
    .ZN(_08525_));
 NOR2_X2 _18182_ (.A1(_08525_),
    .A2(_08507_),
    .ZN(_08526_));
 AND2_X1 _18183_ (.A1(_08506_),
    .A2(_08526_),
    .ZN(_08527_));
 INV_X1 _18184_ (.A(_08527_),
    .ZN(_08528_));
 INV_X1 _18185_ (.A(_08513_),
    .ZN(_08529_));
 OAI221_X1 _18186_ (.A(_08514_),
    .B1(_08520_),
    .B2(_08524_),
    .C1(_08528_),
    .C2(_08529_),
    .ZN(_08530_));
 NOR3_X2 _18187_ (.A1(_08526_),
    .A2(_08504_),
    .A3(_16705_),
    .ZN(_08531_));
 INV_X1 _18188_ (.A(_16704_),
    .ZN(_08532_));
 NOR2_X1 _18189_ (.A1(_08532_),
    .A2(_16703_),
    .ZN(_08533_));
 BUF_X2 _18190_ (.A(_08533_),
    .Z(_08534_));
 INV_X1 _18191_ (.A(_08534_),
    .ZN(_08535_));
 AND2_X1 _18192_ (.A1(_08531_),
    .A2(_08535_),
    .ZN(_08536_));
 INV_X1 _18193_ (.A(_16707_),
    .ZN(_08537_));
 NOR2_X1 _18194_ (.A1(_08537_),
    .A2(_16708_),
    .ZN(_08538_));
 CLKBUF_X2 _18195_ (.A(_08538_),
    .Z(_08539_));
 NOR2_X2 _18196_ (.A1(_16710_),
    .A2(_16709_),
    .ZN(_08540_));
 AND2_X2 _18197_ (.A1(_08539_),
    .A2(_08540_),
    .ZN(_08541_));
 BUF_X2 _18198_ (.A(_08541_),
    .Z(_08542_));
 AND2_X1 _18199_ (.A1(_08536_),
    .A2(_08542_),
    .ZN(_08543_));
 AND2_X1 _18200_ (.A1(_08516_),
    .A2(_16703_),
    .ZN(_08544_));
 INV_X1 _18201_ (.A(_16709_),
    .ZN(_08545_));
 NOR2_X1 _18202_ (.A1(_08545_),
    .A2(_16710_),
    .ZN(_08546_));
 AND2_X1 _18203_ (.A1(_08546_),
    .A2(_08521_),
    .ZN(_08547_));
 CLKBUF_X2 _18204_ (.A(_08547_),
    .Z(_08548_));
 BUF_X2 _18205_ (.A(_08548_),
    .Z(_08549_));
 NAND2_X1 _18206_ (.A1(_08544_),
    .A2(_08549_),
    .ZN(_08550_));
 NOR2_X2 _18207_ (.A1(_16706_),
    .A2(_16705_),
    .ZN(_08551_));
 AND2_X1 _18208_ (.A1(_08508_),
    .A2(_08551_),
    .ZN(_08552_));
 BUF_X2 _18209_ (.A(_08552_),
    .Z(_08553_));
 NAND2_X1 _18210_ (.A1(_08548_),
    .A2(_08553_),
    .ZN(_08554_));
 NAND2_X1 _18211_ (.A1(_08550_),
    .A2(_08554_),
    .ZN(_08555_));
 AND2_X1 _18212_ (.A1(_08551_),
    .A2(_08532_),
    .ZN(_08556_));
 INV_X1 _18213_ (.A(_08556_),
    .ZN(_08557_));
 INV_X1 _18214_ (.A(_08548_),
    .ZN(_08558_));
 AND2_X1 _18215_ (.A1(_08546_),
    .A2(_08512_),
    .ZN(_08559_));
 INV_X1 _18216_ (.A(_08559_),
    .ZN(_08560_));
 AOI21_X1 _18217_ (.A(_08557_),
    .B1(_08558_),
    .B2(_08560_),
    .ZN(_08561_));
 NOR4_X1 _18218_ (.A1(_08530_),
    .A2(_08543_),
    .A3(_08555_),
    .A4(_08561_),
    .ZN(_08562_));
 AND2_X1 _18219_ (.A1(_08537_),
    .A2(_16708_),
    .ZN(_08563_));
 AND2_X1 _18220_ (.A1(_08563_),
    .A2(_08546_),
    .ZN(_08564_));
 BUF_X2 _18221_ (.A(_08564_),
    .Z(_08565_));
 AND2_X1 _18222_ (.A1(_16706_),
    .A2(_16705_),
    .ZN(_08566_));
 CLKBUF_X2 _18223_ (.A(_08566_),
    .Z(_08567_));
 AND2_X2 _18224_ (.A1(_08534_),
    .A2(_08567_),
    .ZN(_08568_));
 NAND2_X1 _18225_ (.A1(_08565_),
    .A2(_08568_),
    .ZN(_08569_));
 AND2_X1 _18226_ (.A1(_08545_),
    .A2(_16710_),
    .ZN(_08570_));
 AND2_X1 _18227_ (.A1(_08563_),
    .A2(_08570_),
    .ZN(_08571_));
 CLKBUF_X2 _18228_ (.A(_08571_),
    .Z(_08572_));
 AND2_X2 _18229_ (.A1(_08509_),
    .A2(_08567_),
    .ZN(_08573_));
 BUF_X2 _18230_ (.A(_08532_),
    .Z(_08574_));
 AND2_X1 _18231_ (.A1(_08567_),
    .A2(_08574_),
    .ZN(_08575_));
 OAI21_X1 _18232_ (.A(_08572_),
    .B1(_08573_),
    .B2(_08575_),
    .ZN(_08576_));
 AND2_X1 _18233_ (.A1(_08506_),
    .A2(_08532_),
    .ZN(_08577_));
 BUF_X2 _18234_ (.A(_08577_),
    .Z(_08578_));
 CLKBUF_X2 _18235_ (.A(_16703_),
    .Z(_08579_));
 CLKBUF_X2 _18236_ (.A(_08570_),
    .Z(_08580_));
 CLKBUF_X2 _18237_ (.A(_08563_),
    .Z(_08581_));
 NAND4_X1 _18238_ (.A1(_08578_),
    .A2(_08579_),
    .A3(_08580_),
    .A4(_08581_),
    .ZN(_08582_));
 AND2_X1 _18239_ (.A1(_08576_),
    .A2(_08582_),
    .ZN(_08583_));
 AND2_X1 _18240_ (.A1(_08563_),
    .A2(_08540_),
    .ZN(_08584_));
 CLKBUF_X2 _18241_ (.A(_08584_),
    .Z(_08585_));
 BUF_X2 _18242_ (.A(_08585_),
    .Z(_08586_));
 INV_X1 _18243_ (.A(_08518_),
    .ZN(_08587_));
 AND2_X1 _18244_ (.A1(_08587_),
    .A2(_08517_),
    .ZN(_08588_));
 INV_X1 _18245_ (.A(_08508_),
    .ZN(_08589_));
 CLKBUF_X2 _18246_ (.A(_08589_),
    .Z(_08590_));
 NAND3_X1 _18247_ (.A1(_08586_),
    .A2(_08588_),
    .A3(_08590_),
    .ZN(_08591_));
 BUF_X2 _18248_ (.A(_08513_),
    .Z(_08592_));
 CLKBUF_X2 _18249_ (.A(_08551_),
    .Z(_08593_));
 AND2_X2 _18250_ (.A1(_08534_),
    .A2(_08593_),
    .ZN(_08594_));
 NOR3_X1 _18251_ (.A1(_08509_),
    .A2(_08504_),
    .A3(_08515_),
    .ZN(_08595_));
 OAI21_X1 _18252_ (.A(_08592_),
    .B1(_08594_),
    .B2(_08595_),
    .ZN(_08596_));
 AND4_X1 _18253_ (.A1(_08569_),
    .A2(_08583_),
    .A3(_08591_),
    .A4(_08596_),
    .ZN(_08597_));
 AND2_X1 _18254_ (.A1(_08540_),
    .A2(_08512_),
    .ZN(_08598_));
 CLKBUF_X2 _18255_ (.A(_08598_),
    .Z(_08599_));
 AND2_X1 _18256_ (.A1(_08551_),
    .A2(_08507_),
    .ZN(_08600_));
 CLKBUF_X2 _18257_ (.A(_08600_),
    .Z(_08601_));
 AND2_X1 _18258_ (.A1(_08599_),
    .A2(_08601_),
    .ZN(_08602_));
 AOI21_X1 _18259_ (.A(_08602_),
    .B1(_08573_),
    .B2(_08585_),
    .ZN(_08603_));
 AND2_X1 _18260_ (.A1(_08580_),
    .A2(_08538_),
    .ZN(_08604_));
 BUF_X2 _18261_ (.A(_08604_),
    .Z(_08605_));
 AND2_X2 _18262_ (.A1(_08567_),
    .A2(_08507_),
    .ZN(_08606_));
 BUF_X2 _18263_ (.A(_08606_),
    .Z(_08607_));
 AND2_X1 _18264_ (.A1(_08570_),
    .A2(_08521_),
    .ZN(_08608_));
 BUF_X2 _18265_ (.A(_08608_),
    .Z(_08609_));
 INV_X1 _18266_ (.A(_08551_),
    .ZN(_08610_));
 NOR2_X1 _18267_ (.A1(_08610_),
    .A2(_08526_),
    .ZN(_08611_));
 AOI22_X1 _18268_ (.A1(_08605_),
    .A2(_08607_),
    .B1(_08609_),
    .B2(_08611_),
    .ZN(_08612_));
 AND2_X1 _18269_ (.A1(_08551_),
    .A2(_16703_),
    .ZN(_08613_));
 BUF_X2 _18270_ (.A(_08517_),
    .Z(_08614_));
 BUF_X2 _18271_ (.A(_08614_),
    .Z(_08615_));
 OAI21_X1 _18272_ (.A(_08565_),
    .B1(_08613_),
    .B2(_08615_),
    .ZN(_08616_));
 INV_X1 _18273_ (.A(_08506_),
    .ZN(_08617_));
 CLKBUF_X2 _18274_ (.A(_08534_),
    .Z(_08618_));
 NOR2_X1 _18275_ (.A1(_08617_),
    .A2(_08618_),
    .ZN(_08619_));
 AND2_X1 _18276_ (.A1(_08516_),
    .A2(_08507_),
    .ZN(_08620_));
 BUF_X2 _18277_ (.A(_08620_),
    .Z(_08621_));
 BUF_X2 _18278_ (.A(_08598_),
    .Z(_08622_));
 AOI22_X1 _18279_ (.A1(_08619_),
    .A2(_08565_),
    .B1(_08621_),
    .B2(_08622_),
    .ZN(_08623_));
 AND4_X1 _18280_ (.A1(_08603_),
    .A2(_08612_),
    .A3(_08616_),
    .A4(_08623_),
    .ZN(_08624_));
 AND2_X1 _18281_ (.A1(_08521_),
    .A2(_08540_),
    .ZN(_08625_));
 AND2_X1 _18282_ (.A1(_08594_),
    .A2(_08625_),
    .ZN(_08626_));
 AND2_X1 _18283_ (.A1(_08625_),
    .A2(_08613_),
    .ZN(_08627_));
 NOR2_X1 _18284_ (.A1(_08626_),
    .A2(_08627_),
    .ZN(_08628_));
 BUF_X2 _18285_ (.A(_08559_),
    .Z(_08629_));
 OAI21_X1 _18286_ (.A(_08629_),
    .B1(_08568_),
    .B2(_08575_),
    .ZN(_08630_));
 CLKBUF_X2 _18287_ (.A(_08506_),
    .Z(_08631_));
 CLKBUF_X2 _18288_ (.A(_08546_),
    .Z(_08632_));
 BUF_X2 _18289_ (.A(_08512_),
    .Z(_08633_));
 NAND4_X1 _18290_ (.A1(_08631_),
    .A2(_08632_),
    .A3(_08579_),
    .A4(_08633_),
    .ZN(_08634_));
 AND2_X1 _18291_ (.A1(_08630_),
    .A2(_08634_),
    .ZN(_08635_));
 BUF_X2 _18292_ (.A(_08625_),
    .Z(_08636_));
 BUF_X2 _18293_ (.A(_08567_),
    .Z(_08637_));
 NAND3_X1 _18294_ (.A1(_08636_),
    .A2(_08535_),
    .A3(_08637_),
    .ZN(_08638_));
 AND2_X1 _18295_ (.A1(_08566_),
    .A2(_08518_),
    .ZN(_08639_));
 CLKBUF_X2 _18296_ (.A(_08639_),
    .Z(_08640_));
 BUF_X2 _18297_ (.A(_08580_),
    .Z(_08641_));
 BUF_X2 _18298_ (.A(_08521_),
    .Z(_08642_));
 NAND3_X1 _18299_ (.A1(_08640_),
    .A2(_08641_),
    .A3(_08642_),
    .ZN(_08643_));
 AND4_X1 _18300_ (.A1(_08628_),
    .A2(_08635_),
    .A3(_08638_),
    .A4(_08643_),
    .ZN(_08644_));
 AND4_X1 _18301_ (.A1(_08562_),
    .A2(_08597_),
    .A3(_08624_),
    .A4(_08644_),
    .ZN(_08645_));
 BUF_X2 _18302_ (.A(_08523_),
    .Z(_08646_));
 AOI21_X1 _18303_ (.A(_08504_),
    .B1(_08535_),
    .B2(_16705_),
    .ZN(_08647_));
 OAI21_X1 _18304_ (.A(_08646_),
    .B1(_08647_),
    .B2(_08601_),
    .ZN(_08648_));
 AND2_X1 _18305_ (.A1(_08580_),
    .A2(_08512_),
    .ZN(_08649_));
 BUF_X2 _18306_ (.A(_08649_),
    .Z(_08650_));
 CLKBUF_X2 _18307_ (.A(_08525_),
    .Z(_08651_));
 INV_X1 _18308_ (.A(_08567_),
    .ZN(_08652_));
 CLKBUF_X2 _18309_ (.A(_08518_),
    .Z(_08653_));
 OAI22_X1 _18310_ (.A1(_08617_),
    .A2(_08651_),
    .B1(_08652_),
    .B2(_08653_),
    .ZN(_08654_));
 AND2_X1 _18311_ (.A1(_08593_),
    .A2(_08651_),
    .ZN(_08655_));
 OAI21_X1 _18312_ (.A(_08650_),
    .B1(_08654_),
    .B2(_08655_),
    .ZN(_08656_));
 CLKBUF_X2 _18313_ (.A(_08540_),
    .Z(_08657_));
 NAND3_X1 _18314_ (.A1(_08601_),
    .A2(_08657_),
    .A3(_08539_),
    .ZN(_08658_));
 NAND3_X1 _18315_ (.A1(_08588_),
    .A2(_08542_),
    .A3(_08590_),
    .ZN(_08659_));
 AND4_X1 _18316_ (.A1(_08648_),
    .A2(_08656_),
    .A3(_08658_),
    .A4(_08659_),
    .ZN(_08660_));
 AND2_X1 _18317_ (.A1(_08567_),
    .A2(_08525_),
    .ZN(_08661_));
 AND2_X1 _18318_ (.A1(_08538_),
    .A2(_08546_),
    .ZN(_08662_));
 CLKBUF_X2 _18319_ (.A(_08662_),
    .Z(_08663_));
 BUF_X2 _18320_ (.A(_08663_),
    .Z(_08664_));
 NOR2_X2 _18321_ (.A1(_08610_),
    .A2(_08533_),
    .ZN(_08665_));
 AOI22_X1 _18322_ (.A1(_08586_),
    .A2(_08661_),
    .B1(_08664_),
    .B2(_08665_),
    .ZN(_08666_));
 AND2_X1 _18323_ (.A1(_08587_),
    .A2(_08505_),
    .ZN(_08667_));
 AOI22_X1 _18324_ (.A1(_08519_),
    .A2(_08572_),
    .B1(_08586_),
    .B2(_08667_),
    .ZN(_08668_));
 INV_X1 _18325_ (.A(_08516_),
    .ZN(_08669_));
 NOR2_X1 _18326_ (.A1(_08669_),
    .A2(_08534_),
    .ZN(_08670_));
 AOI22_X1 _18327_ (.A1(_08609_),
    .A2(_08670_),
    .B1(_08519_),
    .B2(_08629_),
    .ZN(_08671_));
 NOR2_X2 _18328_ (.A1(_08610_),
    .A2(_08509_),
    .ZN(_08672_));
 AOI22_X1 _18329_ (.A1(_08672_),
    .A2(_08586_),
    .B1(_08664_),
    .B2(_08621_),
    .ZN(_08673_));
 AND4_X1 _18330_ (.A1(_08666_),
    .A2(_08668_),
    .A3(_08671_),
    .A4(_08673_),
    .ZN(_08674_));
 CLKBUF_X2 _18331_ (.A(_08511_),
    .Z(_08675_));
 AND2_X2 _18332_ (.A1(_08563_),
    .A2(_08675_),
    .ZN(_08676_));
 BUF_X2 _18333_ (.A(_08676_),
    .Z(_08677_));
 INV_X1 _18334_ (.A(_08552_),
    .ZN(_08678_));
 AND2_X1 _18335_ (.A1(_08518_),
    .A2(_08551_),
    .ZN(_08679_));
 INV_X1 _18336_ (.A(_08679_),
    .ZN(_08680_));
 NAND2_X1 _18337_ (.A1(_08678_),
    .A2(_08680_),
    .ZN(_08681_));
 AND2_X1 _18338_ (.A1(_08567_),
    .A2(_08579_),
    .ZN(_08682_));
 OAI21_X1 _18339_ (.A(_08677_),
    .B1(_08681_),
    .B2(_08682_),
    .ZN(_08683_));
 AND2_X2 _18340_ (.A1(_08516_),
    .A2(_08532_),
    .ZN(_08684_));
 BUF_X2 _18341_ (.A(_08684_),
    .Z(_08685_));
 OAI21_X1 _18342_ (.A(_08677_),
    .B1(_08531_),
    .B2(_08685_),
    .ZN(_08686_));
 NAND2_X1 _18343_ (.A1(_08670_),
    .A2(_08649_),
    .ZN(_08687_));
 AND2_X1 _18344_ (.A1(_08526_),
    .A2(_08551_),
    .ZN(_08688_));
 BUF_X2 _18345_ (.A(_08688_),
    .Z(_08689_));
 NAND2_X1 _18346_ (.A1(_08689_),
    .A2(_08646_),
    .ZN(_08690_));
 AND4_X1 _18347_ (.A1(_08683_),
    .A2(_08686_),
    .A3(_08687_),
    .A4(_08690_),
    .ZN(_08691_));
 NAND4_X2 _18348_ (.A1(_08645_),
    .A2(_08660_),
    .A3(_08674_),
    .A4(_08691_),
    .ZN(_08692_));
 INV_X1 _18349_ (.A(_08510_),
    .ZN(_08693_));
 INV_X1 _18350_ (.A(_08568_),
    .ZN(_08694_));
 AOI21_X1 _18351_ (.A(_08558_),
    .B1(_08693_),
    .B2(_08694_),
    .ZN(_08695_));
 AND2_X2 _18352_ (.A1(_08622_),
    .A2(_08679_),
    .ZN(_08696_));
 AND2_X1 _18353_ (.A1(_08526_),
    .A2(_08567_),
    .ZN(_08697_));
 BUF_X2 _18354_ (.A(_08697_),
    .Z(_08698_));
 AND2_X1 _18355_ (.A1(_08698_),
    .A2(_08549_),
    .ZN(_08699_));
 NOR3_X1 _18356_ (.A1(_08695_),
    .A2(_08696_),
    .A3(_08699_),
    .ZN(_08700_));
 AND2_X1 _18357_ (.A1(_08539_),
    .A2(_08511_),
    .ZN(_08701_));
 BUF_X2 _18358_ (.A(_08701_),
    .Z(_08702_));
 BUF_X2 _18359_ (.A(_08702_),
    .Z(_08703_));
 AND2_X2 _18360_ (.A1(_08526_),
    .A2(_08517_),
    .ZN(_08704_));
 OR3_X1 _18361_ (.A1(_08697_),
    .A2(_08704_),
    .A3(_08594_),
    .ZN(_08705_));
 OAI21_X1 _18362_ (.A(_08703_),
    .B1(_08705_),
    .B2(_08647_),
    .ZN(_08706_));
 AND2_X1 _18363_ (.A1(_08506_),
    .A2(_08507_),
    .ZN(_08707_));
 BUF_X2 _18364_ (.A(_08707_),
    .Z(_08708_));
 NOR2_X1 _18365_ (.A1(_08708_),
    .A2(_08568_),
    .ZN(_08709_));
 INV_X1 _18366_ (.A(_08697_),
    .ZN(_08710_));
 INV_X1 _18367_ (.A(_08704_),
    .ZN(_08711_));
 NAND4_X1 _18368_ (.A1(_08709_),
    .A2(_08710_),
    .A3(_08711_),
    .A4(_08528_),
    .ZN(_08712_));
 NAND2_X1 _18369_ (.A1(_08712_),
    .A2(_08622_),
    .ZN(_08713_));
 AND2_X2 _18370_ (.A1(_08534_),
    .A2(_08517_),
    .ZN(_08714_));
 AND2_X1 _18371_ (.A1(_08506_),
    .A2(_08653_),
    .ZN(_08715_));
 OAI21_X1 _18372_ (.A(_08636_),
    .B1(_08714_),
    .B2(_08715_),
    .ZN(_08716_));
 NAND3_X1 _18373_ (.A1(_08605_),
    .A2(_08672_),
    .A3(_08587_),
    .ZN(_08717_));
 AND2_X1 _18374_ (.A1(_08506_),
    .A2(_16703_),
    .ZN(_08718_));
 OAI21_X1 _18375_ (.A(_08664_),
    .B1(_08718_),
    .B2(_08573_),
    .ZN(_08719_));
 AND3_X1 _18376_ (.A1(_08716_),
    .A2(_08717_),
    .A3(_08719_),
    .ZN(_08720_));
 NAND4_X2 _18377_ (.A1(_08700_),
    .A2(_08706_),
    .A3(_08713_),
    .A4(_08720_),
    .ZN(_08721_));
 NOR2_X2 _18378_ (.A1(_08692_),
    .A2(_08721_),
    .ZN(_08722_));
 OAI21_X1 _18379_ (.A(_08646_),
    .B1(_08527_),
    .B2(_08661_),
    .ZN(_08723_));
 CLKBUF_X2 _18380_ (.A(_08556_),
    .Z(_08724_));
 AND2_X1 _18381_ (.A1(_08676_),
    .A2(_08724_),
    .ZN(_08725_));
 NAND3_X1 _18382_ (.A1(_08620_),
    .A2(_08675_),
    .A3(_08563_),
    .ZN(_08726_));
 INV_X1 _18383_ (.A(_08676_),
    .ZN(_08727_));
 OAI21_X1 _18384_ (.A(_08726_),
    .B1(_08727_),
    .B2(_08711_),
    .ZN(_08728_));
 AOI211_X1 _18385_ (.A(_08725_),
    .B(_08728_),
    .C1(_08594_),
    .C2(_08676_),
    .ZN(_08729_));
 OAI21_X1 _18386_ (.A(_08523_),
    .B1(_08685_),
    .B2(_08672_),
    .ZN(_08730_));
 INV_X1 _18387_ (.A(_08526_),
    .ZN(_08731_));
 NOR2_X2 _18388_ (.A1(_08652_),
    .A2(_08534_),
    .ZN(_08732_));
 BUF_X2 _18389_ (.A(_08631_),
    .Z(_08733_));
 OAI211_X1 _18390_ (.A(_08676_),
    .B(_08731_),
    .C1(_08732_),
    .C2(_08733_),
    .ZN(_08734_));
 AND4_X1 _18391_ (.A1(_08723_),
    .A2(_08729_),
    .A3(_08730_),
    .A4(_08734_),
    .ZN(_08735_));
 OAI21_X1 _18392_ (.A(_08592_),
    .B1(_08588_),
    .B2(_08679_),
    .ZN(_08736_));
 AND2_X1 _18393_ (.A1(_08606_),
    .A2(_08513_),
    .ZN(_08737_));
 AND2_X1 _18394_ (.A1(_08577_),
    .A2(_08513_),
    .ZN(_08738_));
 AOI211_X1 _18395_ (.A(_08737_),
    .B(_08738_),
    .C1(_08698_),
    .C2(_08592_),
    .ZN(_08739_));
 OAI21_X1 _18396_ (.A(_08703_),
    .B1(_08732_),
    .B2(_08510_),
    .ZN(_08740_));
 NAND2_X1 _18397_ (.A1(_08594_),
    .A2(_08702_),
    .ZN(_08741_));
 NAND2_X1 _18398_ (.A1(_08714_),
    .A2(_08702_),
    .ZN(_08742_));
 AND2_X1 _18399_ (.A1(_08741_),
    .A2(_08742_),
    .ZN(_08743_));
 AND4_X1 _18400_ (.A1(_08736_),
    .A2(_08739_),
    .A3(_08740_),
    .A4(_08743_),
    .ZN(_08744_));
 OAI21_X1 _18401_ (.A(_08605_),
    .B1(_08621_),
    .B2(_08613_),
    .ZN(_08745_));
 AND2_X1 _18402_ (.A1(_08667_),
    .A2(_08589_),
    .ZN(_08746_));
 OR2_X1 _18403_ (.A1(_08573_),
    .A2(_08639_),
    .ZN(_08747_));
 OAI21_X1 _18404_ (.A(_08605_),
    .B1(_08746_),
    .B2(_08747_),
    .ZN(_08748_));
 NAND3_X1 _18405_ (.A1(_08578_),
    .A2(_08633_),
    .A3(_08641_),
    .ZN(_08749_));
 OAI21_X1 _18406_ (.A(_08650_),
    .B1(_08681_),
    .B2(_08704_),
    .ZN(_08750_));
 AND4_X1 _18407_ (.A1(_08745_),
    .A2(_08748_),
    .A3(_08749_),
    .A4(_08750_),
    .ZN(_08751_));
 INV_X1 _18408_ (.A(_08571_),
    .ZN(_08752_));
 AOI221_X4 _18409_ (.A(_08752_),
    .B1(_08507_),
    .B2(_08535_),
    .C1(_08617_),
    .C2(_08652_),
    .ZN(_08753_));
 INV_X1 _18410_ (.A(_08608_),
    .ZN(_08754_));
 NOR2_X1 _18411_ (.A1(_08709_),
    .A2(_08754_),
    .ZN(_08755_));
 AND2_X1 _18412_ (.A1(_08571_),
    .A2(_08679_),
    .ZN(_08756_));
 NAND2_X1 _18413_ (.A1(_08609_),
    .A2(_08684_),
    .ZN(_08757_));
 AND2_X2 _18414_ (.A1(_08517_),
    .A2(_08509_),
    .ZN(_08758_));
 NAND2_X1 _18415_ (.A1(_08609_),
    .A2(_08758_),
    .ZN(_08759_));
 OAI211_X1 _18416_ (.A(_08757_),
    .B(_08759_),
    .C1(_08754_),
    .C2(_08557_),
    .ZN(_08760_));
 NOR4_X1 _18417_ (.A1(_08753_),
    .A2(_08755_),
    .A3(_08756_),
    .A4(_08760_),
    .ZN(_08761_));
 NAND4_X2 _18418_ (.A1(_08735_),
    .A2(_08744_),
    .A3(_08751_),
    .A4(_08761_),
    .ZN(_08762_));
 AND2_X1 _18419_ (.A1(_08578_),
    .A2(_08548_),
    .ZN(_08763_));
 AND2_X1 _18420_ (.A1(_08506_),
    .A2(_08534_),
    .ZN(_08764_));
 AND2_X1 _18421_ (.A1(_08764_),
    .A2(_08548_),
    .ZN(_08765_));
 NOR2_X1 _18422_ (.A1(_08763_),
    .A2(_08765_),
    .ZN(_08766_));
 INV_X1 _18423_ (.A(_08564_),
    .ZN(_08767_));
 INV_X1 _18424_ (.A(_08606_),
    .ZN(_08768_));
 AOI21_X1 _18425_ (.A(_08767_),
    .B1(_08528_),
    .B2(_08768_),
    .ZN(_08769_));
 AND2_X1 _18426_ (.A1(_08564_),
    .A2(_08601_),
    .ZN(_08770_));
 AND2_X1 _18427_ (.A1(_08564_),
    .A2(_08758_),
    .ZN(_08771_));
 AND2_X1 _18428_ (.A1(_08564_),
    .A2(_08556_),
    .ZN(_08772_));
 NOR4_X1 _18429_ (.A1(_08769_),
    .A2(_08770_),
    .A3(_08771_),
    .A4(_08772_),
    .ZN(_08773_));
 NOR2_X1 _18430_ (.A1(_08652_),
    .A2(_08653_),
    .ZN(_08774_));
 AND2_X1 _18431_ (.A1(_08774_),
    .A2(_08548_),
    .ZN(_08775_));
 INV_X1 _18432_ (.A(_08775_),
    .ZN(_08776_));
 AND2_X1 _18433_ (.A1(_08547_),
    .A2(_08613_),
    .ZN(_08777_));
 AND2_X1 _18434_ (.A1(_08758_),
    .A2(_08548_),
    .ZN(_08778_));
 AOI211_X1 _18435_ (.A(_08777_),
    .B(_08778_),
    .C1(_08685_),
    .C2(_08548_),
    .ZN(_08779_));
 AND4_X1 _18436_ (.A1(_08766_),
    .A2(_08773_),
    .A3(_08776_),
    .A4(_08779_),
    .ZN(_08780_));
 AND2_X1 _18437_ (.A1(_08704_),
    .A2(_08663_),
    .ZN(_08781_));
 AND2_X1 _18438_ (.A1(_08714_),
    .A2(_08663_),
    .ZN(_08782_));
 AOI211_X1 _18439_ (.A(_08781_),
    .B(_08782_),
    .C1(_08663_),
    .C2(_08613_),
    .ZN(_08783_));
 OAI21_X1 _18440_ (.A(_08663_),
    .B1(_08746_),
    .B2(_08573_),
    .ZN(_08784_));
 OAI21_X1 _18441_ (.A(_08629_),
    .B1(_08689_),
    .B2(_08758_),
    .ZN(_08785_));
 OAI21_X1 _18442_ (.A(_08629_),
    .B1(_08708_),
    .B2(_08682_),
    .ZN(_08786_));
 AND4_X1 _18443_ (.A1(_08783_),
    .A2(_08784_),
    .A3(_08785_),
    .A4(_08786_),
    .ZN(_08787_));
 AND3_X1 _18444_ (.A1(_08670_),
    .A2(_08731_),
    .A3(_08541_),
    .ZN(_08788_));
 INV_X1 _18445_ (.A(_08788_),
    .ZN(_08789_));
 NAND3_X1 _18446_ (.A1(_08724_),
    .A2(_08657_),
    .A3(_08539_),
    .ZN(_08790_));
 NAND4_X1 _18447_ (.A1(_08618_),
    .A2(_08539_),
    .A3(_08657_),
    .A4(_08593_),
    .ZN(_08791_));
 NAND3_X1 _18448_ (.A1(_08789_),
    .A2(_08790_),
    .A3(_08791_),
    .ZN(_08792_));
 INV_X1 _18449_ (.A(_08541_),
    .ZN(_08793_));
 BUF_X2 _18450_ (.A(_08507_),
    .Z(_08794_));
 AOI211_X1 _18451_ (.A(_08652_),
    .B(_08793_),
    .C1(_08651_),
    .C2(_08794_),
    .ZN(_08795_));
 NAND4_X1 _18452_ (.A1(_08599_),
    .A2(_08535_),
    .A3(_08731_),
    .A4(_08614_),
    .ZN(_08796_));
 BUF_X2 _18453_ (.A(_08575_),
    .Z(_08797_));
 NAND2_X1 _18454_ (.A1(_08797_),
    .A2(_08599_),
    .ZN(_08798_));
 NAND3_X1 _18455_ (.A1(_08599_),
    .A2(_08618_),
    .A3(_08637_),
    .ZN(_08799_));
 NAND3_X1 _18456_ (.A1(_08796_),
    .A2(_08798_),
    .A3(_08799_),
    .ZN(_08800_));
 INV_X1 _18457_ (.A(_08707_),
    .ZN(_08801_));
 INV_X2 _18458_ (.A(_08578_),
    .ZN(_08802_));
 AOI21_X1 _18459_ (.A(_08793_),
    .B1(_08801_),
    .B2(_08802_),
    .ZN(_08803_));
 NOR4_X1 _18460_ (.A1(_08792_),
    .A2(_08795_),
    .A3(_08800_),
    .A4(_08803_),
    .ZN(_08804_));
 OAI21_X1 _18461_ (.A(_08636_),
    .B1(_08708_),
    .B2(_08661_),
    .ZN(_08805_));
 OAI21_X1 _18462_ (.A(_08585_),
    .B1(_08667_),
    .B2(_08698_),
    .ZN(_08806_));
 OAI21_X1 _18463_ (.A(_08585_),
    .B1(_08621_),
    .B2(_08672_),
    .ZN(_08807_));
 OAI211_X1 _18464_ (.A(_08636_),
    .B(_08579_),
    .C1(_08615_),
    .C2(_08593_),
    .ZN(_08808_));
 AND4_X1 _18465_ (.A1(_08805_),
    .A2(_08806_),
    .A3(_08807_),
    .A4(_08808_),
    .ZN(_08809_));
 NAND4_X2 _18466_ (.A1(_08780_),
    .A2(_08787_),
    .A3(_08804_),
    .A4(_08809_),
    .ZN(_08810_));
 NOR2_X2 _18467_ (.A1(_08762_),
    .A2(_08810_),
    .ZN(_08811_));
 NAND2_X1 _18468_ (.A1(_08722_),
    .A2(_08811_),
    .ZN(_08812_));
 OAI22_X1 _18469_ (.A1(_08692_),
    .A2(_08721_),
    .B1(_08762_),
    .B2(_08810_),
    .ZN(_08813_));
 NAND2_X1 _18470_ (.A1(_08812_),
    .A2(_08813_),
    .ZN(_08814_));
 XNOR2_X1 _18471_ (.A(_08503_),
    .B(_08814_),
    .ZN(_08815_));
 INV_X1 _18472_ (.A(_16793_),
    .ZN(_08816_));
 NOR2_X1 _18473_ (.A1(_08816_),
    .A2(_16794_),
    .ZN(_08817_));
 INV_X1 _18474_ (.A(_08817_),
    .ZN(_08818_));
 INV_X1 _18475_ (.A(_16792_),
    .ZN(_08819_));
 NOR2_X2 _18476_ (.A1(_08819_),
    .A2(_16791_),
    .ZN(_08820_));
 NOR2_X2 _18477_ (.A1(_08818_),
    .A2(_08820_),
    .ZN(_08821_));
 INV_X1 _18478_ (.A(_16791_),
    .ZN(_08822_));
 NOR2_X2 _18479_ (.A1(_08822_),
    .A2(_16792_),
    .ZN(_08823_));
 INV_X2 _18480_ (.A(_08823_),
    .ZN(_08824_));
 NOR2_X2 _18481_ (.A1(_16798_),
    .A2(_16797_),
    .ZN(_08825_));
 NOR2_X1 _18482_ (.A1(_16796_),
    .A2(_16795_),
    .ZN(_08826_));
 CLKBUF_X2 _18483_ (.A(_08826_),
    .Z(_08827_));
 AND2_X1 _18484_ (.A1(_08825_),
    .A2(_08827_),
    .ZN(_08828_));
 BUF_X2 _18485_ (.A(_08828_),
    .Z(_08829_));
 BUF_X2 _18486_ (.A(_08829_),
    .Z(_08830_));
 NAND3_X1 _18487_ (.A1(_08821_),
    .A2(_08824_),
    .A3(_08830_),
    .ZN(_08831_));
 INV_X1 _18488_ (.A(_16795_),
    .ZN(_08832_));
 NOR2_X2 _18489_ (.A1(_08832_),
    .A2(_16796_),
    .ZN(_08833_));
 AND2_X2 _18490_ (.A1(_08833_),
    .A2(_08825_),
    .ZN(_08834_));
 NOR2_X2 _18491_ (.A1(_16794_),
    .A2(_16793_),
    .ZN(_08835_));
 AND2_X1 _18492_ (.A1(_08835_),
    .A2(_08819_),
    .ZN(_08836_));
 AND2_X1 _18493_ (.A1(_08834_),
    .A2(_08836_),
    .ZN(_08837_));
 AND2_X2 _18494_ (.A1(_08820_),
    .A2(_08835_),
    .ZN(_08838_));
 AND2_X1 _18495_ (.A1(_08821_),
    .A2(_08834_),
    .ZN(_08839_));
 AOI221_X4 _18496_ (.A(_08837_),
    .B1(_08834_),
    .B2(_08838_),
    .C1(_08839_),
    .C2(_08824_),
    .ZN(_08840_));
 AND2_X1 _18497_ (.A1(_16794_),
    .A2(_16793_),
    .ZN(_08841_));
 CLKBUF_X2 _18498_ (.A(_08841_),
    .Z(_08842_));
 BUF_X2 _18499_ (.A(_08842_),
    .Z(_08843_));
 CLKBUF_X2 _18500_ (.A(_08822_),
    .Z(_08844_));
 CLKBUF_X2 _18501_ (.A(_08819_),
    .Z(_08845_));
 OAI211_X1 _18502_ (.A(_08829_),
    .B(_08843_),
    .C1(_08844_),
    .C2(_08845_),
    .ZN(_08846_));
 CLKBUF_X2 _18503_ (.A(_08834_),
    .Z(_08847_));
 INV_X1 _18504_ (.A(_16794_),
    .ZN(_08848_));
 NOR2_X1 _18505_ (.A1(_08848_),
    .A2(_16793_),
    .ZN(_08849_));
 AND2_X1 _18506_ (.A1(_08849_),
    .A2(_08845_),
    .ZN(_08850_));
 NAND2_X1 _18507_ (.A1(_08847_),
    .A2(_08850_),
    .ZN(_08851_));
 AND2_X1 _18508_ (.A1(_08849_),
    .A2(_16792_),
    .ZN(_08852_));
 CLKBUF_X2 _18509_ (.A(_08852_),
    .Z(_08853_));
 NAND2_X1 _18510_ (.A1(_08847_),
    .A2(_08853_),
    .ZN(_08854_));
 AND2_X2 _18511_ (.A1(_08841_),
    .A2(_08819_),
    .ZN(_08855_));
 NAND2_X1 _18512_ (.A1(_08834_),
    .A2(_08855_),
    .ZN(_08856_));
 AND2_X1 _18513_ (.A1(_16791_),
    .A2(_16792_),
    .ZN(_08857_));
 BUF_X2 _18514_ (.A(_08857_),
    .Z(_08858_));
 AND2_X1 _18515_ (.A1(_08858_),
    .A2(_08842_),
    .ZN(_08859_));
 BUF_X2 _18516_ (.A(_08859_),
    .Z(_08860_));
 NAND2_X1 _18517_ (.A1(_08834_),
    .A2(_08860_),
    .ZN(_08861_));
 AND4_X1 _18518_ (.A1(_08851_),
    .A2(_08854_),
    .A3(_08856_),
    .A4(_08861_),
    .ZN(_08862_));
 AND4_X1 _18519_ (.A1(_08831_),
    .A2(_08840_),
    .A3(_08846_),
    .A4(_08862_),
    .ZN(_08863_));
 AND2_X1 _18520_ (.A1(_08832_),
    .A2(_16796_),
    .ZN(_08864_));
 AND2_X1 _18521_ (.A1(_08864_),
    .A2(_08825_),
    .ZN(_08865_));
 INV_X1 _18522_ (.A(_08865_),
    .ZN(_08866_));
 INV_X2 _18523_ (.A(_08857_),
    .ZN(_08867_));
 BUF_X2 _18524_ (.A(_08835_),
    .Z(_08868_));
 NAND2_X1 _18525_ (.A1(_08867_),
    .A2(_08868_),
    .ZN(_08869_));
 NOR2_X1 _18526_ (.A1(_08866_),
    .A2(_08869_),
    .ZN(_08870_));
 INV_X1 _18527_ (.A(_08870_),
    .ZN(_08871_));
 NOR2_X1 _18528_ (.A1(_16791_),
    .A2(_16792_),
    .ZN(_08872_));
 INV_X1 _18529_ (.A(_08872_),
    .ZN(_08873_));
 CLKBUF_X2 _18530_ (.A(_08849_),
    .Z(_08874_));
 NAND2_X1 _18531_ (.A1(_08873_),
    .A2(_08874_),
    .ZN(_08875_));
 OR2_X1 _18532_ (.A1(_08866_),
    .A2(_08875_),
    .ZN(_08876_));
 CLKBUF_X2 _18533_ (.A(_08817_),
    .Z(_08877_));
 CLKBUF_X2 _18534_ (.A(_16792_),
    .Z(_08878_));
 AND2_X1 _18535_ (.A1(_08877_),
    .A2(_08878_),
    .ZN(_08879_));
 AND2_X1 _18536_ (.A1(_08865_),
    .A2(_08879_),
    .ZN(_08880_));
 INV_X1 _18537_ (.A(_08880_),
    .ZN(_08881_));
 AND2_X2 _18538_ (.A1(_08823_),
    .A2(_08842_),
    .ZN(_08882_));
 NAND2_X1 _18539_ (.A1(_08865_),
    .A2(_08882_),
    .ZN(_08883_));
 NAND4_X1 _18540_ (.A1(_08871_),
    .A2(_08876_),
    .A3(_08881_),
    .A4(_08883_),
    .ZN(_08884_));
 AND2_X1 _18541_ (.A1(_16796_),
    .A2(_16795_),
    .ZN(_08885_));
 CLKBUF_X2 _18542_ (.A(_08885_),
    .Z(_08886_));
 AND2_X1 _18543_ (.A1(_08886_),
    .A2(_08825_),
    .ZN(_08887_));
 BUF_X2 _18544_ (.A(_08887_),
    .Z(_08888_));
 AND2_X2 _18545_ (.A1(_08868_),
    .A2(_16791_),
    .ZN(_08889_));
 AND2_X1 _18546_ (.A1(_08888_),
    .A2(_08889_),
    .ZN(_08890_));
 AND3_X1 _18547_ (.A1(_08887_),
    .A2(_16791_),
    .A3(_08877_),
    .ZN(_08891_));
 INV_X1 _18548_ (.A(_08887_),
    .ZN(_08892_));
 INV_X1 _18549_ (.A(_08853_),
    .ZN(_08893_));
 AND2_X1 _18550_ (.A1(_08842_),
    .A2(_08822_),
    .ZN(_08894_));
 INV_X1 _18551_ (.A(_08894_),
    .ZN(_08895_));
 AOI21_X1 _18552_ (.A(_08892_),
    .B1(_08893_),
    .B2(_08895_),
    .ZN(_08896_));
 NOR4_X1 _18553_ (.A1(_08884_),
    .A2(_08890_),
    .A3(_08891_),
    .A4(_08896_),
    .ZN(_08897_));
 INV_X1 _18554_ (.A(_16798_),
    .ZN(_08898_));
 AND2_X1 _18555_ (.A1(_08898_),
    .A2(_16797_),
    .ZN(_08899_));
 AND2_X1 _18556_ (.A1(_08899_),
    .A2(_08885_),
    .ZN(_08900_));
 CLKBUF_X2 _18557_ (.A(_08900_),
    .Z(_08901_));
 AND2_X1 _18558_ (.A1(_08849_),
    .A2(_08820_),
    .ZN(_08902_));
 CLKBUF_X2 _18559_ (.A(_08902_),
    .Z(_08903_));
 BUF_X2 _18560_ (.A(_08850_),
    .Z(_08904_));
 OAI21_X1 _18561_ (.A(_08901_),
    .B1(_08903_),
    .B2(_08904_),
    .ZN(_08905_));
 AND2_X2 _18562_ (.A1(_08864_),
    .A2(_08899_),
    .ZN(_08906_));
 AND2_X2 _18563_ (.A1(_08874_),
    .A2(_08823_),
    .ZN(_08907_));
 AND2_X1 _18564_ (.A1(_08841_),
    .A2(_16792_),
    .ZN(_08908_));
 BUF_X2 _18565_ (.A(_08908_),
    .Z(_08909_));
 OAI21_X1 _18566_ (.A(_08906_),
    .B1(_08907_),
    .B2(_08909_),
    .ZN(_08910_));
 AND2_X2 _18567_ (.A1(_08877_),
    .A2(_08858_),
    .ZN(_08911_));
 NAND2_X1 _18568_ (.A1(_08906_),
    .A2(_08911_),
    .ZN(_08912_));
 CLKBUF_X2 _18569_ (.A(_08864_),
    .Z(_08913_));
 BUF_X2 _18570_ (.A(_08899_),
    .Z(_08914_));
 AND2_X2 _18571_ (.A1(_08835_),
    .A2(_08878_),
    .ZN(_08915_));
 OAI211_X1 _18572_ (.A(_08913_),
    .B(_08914_),
    .C1(_08836_),
    .C2(_08915_),
    .ZN(_08916_));
 AND3_X1 _18573_ (.A1(_08910_),
    .A2(_08912_),
    .A3(_08916_),
    .ZN(_08917_));
 NAND2_X1 _18574_ (.A1(_08873_),
    .A2(_08841_),
    .ZN(_08918_));
 INV_X1 _18575_ (.A(_08918_),
    .ZN(_08919_));
 AND2_X1 _18576_ (.A1(_08919_),
    .A2(_08901_),
    .ZN(_08920_));
 INV_X1 _18577_ (.A(_08920_),
    .ZN(_08921_));
 NAND2_X1 _18578_ (.A1(_08901_),
    .A2(_08889_),
    .ZN(_08922_));
 AND2_X1 _18579_ (.A1(_08877_),
    .A2(_08845_),
    .ZN(_08923_));
 NAND2_X1 _18580_ (.A1(_08901_),
    .A2(_08923_),
    .ZN(_08924_));
 NAND2_X1 _18581_ (.A1(_08901_),
    .A2(_08911_),
    .ZN(_08925_));
 AND3_X1 _18582_ (.A1(_08922_),
    .A2(_08924_),
    .A3(_08925_),
    .ZN(_08926_));
 AND4_X1 _18583_ (.A1(_08905_),
    .A2(_08917_),
    .A3(_08921_),
    .A4(_08926_),
    .ZN(_08927_));
 AND2_X1 _18584_ (.A1(_08899_),
    .A2(_08833_),
    .ZN(_08928_));
 CLKBUF_X2 _18585_ (.A(_08928_),
    .Z(_08929_));
 AND2_X1 _18586_ (.A1(_08823_),
    .A2(_08877_),
    .ZN(_08930_));
 NAND2_X1 _18587_ (.A1(_08929_),
    .A2(_08930_),
    .ZN(_08931_));
 INV_X1 _18588_ (.A(_08929_),
    .ZN(_08932_));
 AND2_X1 _18589_ (.A1(_08820_),
    .A2(_08817_),
    .ZN(_08933_));
 INV_X1 _18590_ (.A(_08933_),
    .ZN(_08934_));
 OAI21_X1 _18591_ (.A(_08931_),
    .B1(_08932_),
    .B2(_08934_),
    .ZN(_08935_));
 BUF_X2 _18592_ (.A(_08929_),
    .Z(_08936_));
 AOI21_X1 _18593_ (.A(_08935_),
    .B1(_08889_),
    .B2(_08936_),
    .ZN(_08937_));
 NOR2_X2 _18594_ (.A1(_08875_),
    .A2(_08858_),
    .ZN(_08938_));
 OAI21_X1 _18595_ (.A(_08929_),
    .B1(_08938_),
    .B2(_08860_),
    .ZN(_08939_));
 AND2_X1 _18596_ (.A1(_08899_),
    .A2(_08827_),
    .ZN(_08940_));
 BUF_X2 _18597_ (.A(_08940_),
    .Z(_08941_));
 AND2_X1 _18598_ (.A1(_08823_),
    .A2(_08835_),
    .ZN(_08942_));
 BUF_X2 _18599_ (.A(_08942_),
    .Z(_08943_));
 OAI21_X1 _18600_ (.A(_08941_),
    .B1(_08911_),
    .B2(_08943_),
    .ZN(_08944_));
 AND2_X1 _18601_ (.A1(_08842_),
    .A2(_16791_),
    .ZN(_08945_));
 OAI21_X1 _18602_ (.A(_08941_),
    .B1(_08853_),
    .B2(_08945_),
    .ZN(_08946_));
 AND4_X1 _18603_ (.A1(_08937_),
    .A2(_08939_),
    .A3(_08944_),
    .A4(_08946_),
    .ZN(_08947_));
 NAND4_X2 _18604_ (.A1(_08863_),
    .A2(_08897_),
    .A3(_08927_),
    .A4(_08947_),
    .ZN(_08948_));
 AND2_X1 _18605_ (.A1(_16798_),
    .A2(_16797_),
    .ZN(_08949_));
 CLKBUF_X2 _18606_ (.A(_08949_),
    .Z(_08950_));
 AND2_X1 _18607_ (.A1(_08833_),
    .A2(_08950_),
    .ZN(_08951_));
 CLKBUF_X2 _18608_ (.A(_08951_),
    .Z(_08952_));
 NAND2_X1 _18609_ (.A1(_08838_),
    .A2(_08952_),
    .ZN(_08953_));
 CLKBUF_X2 _18610_ (.A(_08933_),
    .Z(_08954_));
 NAND2_X1 _18611_ (.A1(_08954_),
    .A2(_08952_),
    .ZN(_08955_));
 AND2_X1 _18612_ (.A1(_08953_),
    .A2(_08955_),
    .ZN(_08956_));
 AND2_X2 _18613_ (.A1(_08950_),
    .A2(_08826_),
    .ZN(_08957_));
 AND2_X1 _18614_ (.A1(_08882_),
    .A2(_08957_),
    .ZN(_08958_));
 INV_X1 _18615_ (.A(_08958_),
    .ZN(_08959_));
 NAND2_X1 _18616_ (.A1(_08850_),
    .A2(_08957_),
    .ZN(_08960_));
 AND2_X1 _18617_ (.A1(_08957_),
    .A2(_08908_),
    .ZN(_08961_));
 INV_X1 _18618_ (.A(_08961_),
    .ZN(_08962_));
 AND3_X1 _18619_ (.A1(_08877_),
    .A2(_08827_),
    .A3(_08950_),
    .ZN(_08963_));
 CLKBUF_X2 _18620_ (.A(_08872_),
    .Z(_08964_));
 AND2_X1 _18621_ (.A1(_08835_),
    .A2(_08964_),
    .ZN(_08965_));
 AOI22_X1 _18622_ (.A1(_08963_),
    .A2(_08873_),
    .B1(_08957_),
    .B2(_08965_),
    .ZN(_08966_));
 AND4_X1 _18623_ (.A1(_08959_),
    .A2(_08960_),
    .A3(_08962_),
    .A4(_08966_),
    .ZN(_08967_));
 AND2_X1 _18624_ (.A1(_08849_),
    .A2(_08857_),
    .ZN(_08968_));
 CLKBUF_X2 _18625_ (.A(_08968_),
    .Z(_08969_));
 AND2_X1 _18626_ (.A1(_08969_),
    .A2(_08951_),
    .ZN(_08970_));
 INV_X1 _18627_ (.A(_08970_),
    .ZN(_08971_));
 BUF_X2 _18628_ (.A(_08951_),
    .Z(_08972_));
 BUF_X2 _18629_ (.A(_16791_),
    .Z(_08973_));
 OAI211_X1 _18630_ (.A(_08972_),
    .B(_08843_),
    .C1(_08973_),
    .C2(_08845_),
    .ZN(_08974_));
 AND4_X1 _18631_ (.A1(_08956_),
    .A2(_08967_),
    .A3(_08971_),
    .A4(_08974_),
    .ZN(_08975_));
 AND2_X1 _18632_ (.A1(_08864_),
    .A2(_08949_),
    .ZN(_08976_));
 AND2_X1 _18633_ (.A1(_08841_),
    .A2(_08964_),
    .ZN(_08977_));
 AND2_X1 _18634_ (.A1(_08976_),
    .A2(_08977_),
    .ZN(_08978_));
 INV_X1 _18635_ (.A(_08978_),
    .ZN(_08979_));
 AND3_X1 _18636_ (.A1(_08859_),
    .A2(_08913_),
    .A3(_08950_),
    .ZN(_08980_));
 INV_X1 _18637_ (.A(_08980_),
    .ZN(_08981_));
 BUF_X2 _18638_ (.A(_08976_),
    .Z(_08982_));
 INV_X1 _18639_ (.A(_08982_),
    .ZN(_08983_));
 NAND2_X1 _18640_ (.A1(_08824_),
    .A2(_08849_),
    .ZN(_08984_));
 OAI211_X1 _18641_ (.A(_08979_),
    .B(_08981_),
    .C1(_08983_),
    .C2(_08984_),
    .ZN(_08985_));
 BUF_X2 _18642_ (.A(_08930_),
    .Z(_08986_));
 CLKBUF_X2 _18643_ (.A(_08879_),
    .Z(_08987_));
 OAI21_X1 _18644_ (.A(_08982_),
    .B1(_08986_),
    .B2(_08987_),
    .ZN(_08988_));
 BUF_X2 _18645_ (.A(_08836_),
    .Z(_08989_));
 NAND2_X1 _18646_ (.A1(_08982_),
    .A2(_08989_),
    .ZN(_08990_));
 INV_X1 _18647_ (.A(_08838_),
    .ZN(_08991_));
 OAI211_X1 _18648_ (.A(_08988_),
    .B(_08990_),
    .C1(_08983_),
    .C2(_08991_),
    .ZN(_08992_));
 AND2_X1 _18649_ (.A1(_08886_),
    .A2(_08950_),
    .ZN(_08993_));
 CLKBUF_X2 _18650_ (.A(_08993_),
    .Z(_08994_));
 INV_X1 _18651_ (.A(_08994_),
    .ZN(_08995_));
 INV_X1 _18652_ (.A(_08907_),
    .ZN(_08996_));
 AOI21_X1 _18653_ (.A(_08995_),
    .B1(_08996_),
    .B2(_08895_),
    .ZN(_08997_));
 BUF_X2 _18654_ (.A(_08923_),
    .Z(_08998_));
 INV_X1 _18655_ (.A(_08998_),
    .ZN(_08999_));
 AOI21_X1 _18656_ (.A(_08995_),
    .B1(_08999_),
    .B2(_08869_),
    .ZN(_09000_));
 NOR4_X1 _18657_ (.A1(_08985_),
    .A2(_08992_),
    .A3(_08997_),
    .A4(_09000_),
    .ZN(_09001_));
 NOR2_X1 _18658_ (.A1(_08898_),
    .A2(_16797_),
    .ZN(_09002_));
 CLKBUF_X2 _18659_ (.A(_09002_),
    .Z(_09003_));
 AND2_X1 _18660_ (.A1(_09003_),
    .A2(_08827_),
    .ZN(_09004_));
 BUF_X2 _18661_ (.A(_09004_),
    .Z(_09005_));
 NAND2_X1 _18662_ (.A1(_09005_),
    .A2(_08904_),
    .ZN(_09006_));
 AND2_X2 _18663_ (.A1(_08833_),
    .A2(_09003_),
    .ZN(_09007_));
 BUF_X2 _18664_ (.A(_09007_),
    .Z(_09008_));
 BUF_X2 _18665_ (.A(_08977_),
    .Z(_09009_));
 NOR2_X1 _18666_ (.A1(_08860_),
    .A2(_09009_),
    .ZN(_09010_));
 INV_X1 _18667_ (.A(_09010_),
    .ZN(_09011_));
 OAI21_X1 _18668_ (.A(_09008_),
    .B1(_09011_),
    .B2(_08938_),
    .ZN(_09012_));
 OAI21_X1 _18669_ (.A(_09007_),
    .B1(_08987_),
    .B2(_08889_),
    .ZN(_09013_));
 AND2_X1 _18670_ (.A1(_08858_),
    .A2(_08835_),
    .ZN(_09014_));
 INV_X1 _18671_ (.A(_09014_),
    .ZN(_09015_));
 INV_X1 _18672_ (.A(_08965_),
    .ZN(_09016_));
 NAND2_X2 _18673_ (.A1(_09015_),
    .A2(_09016_),
    .ZN(_09017_));
 OAI21_X1 _18674_ (.A(_09005_),
    .B1(_09017_),
    .B2(_08986_),
    .ZN(_09018_));
 AND4_X1 _18675_ (.A1(_09006_),
    .A2(_09012_),
    .A3(_09013_),
    .A4(_09018_),
    .ZN(_09019_));
 AND2_X2 _18676_ (.A1(_09002_),
    .A2(_08885_),
    .ZN(_09020_));
 AND2_X2 _18677_ (.A1(_08820_),
    .A2(_08842_),
    .ZN(_09021_));
 AND2_X1 _18678_ (.A1(_09020_),
    .A2(_09021_),
    .ZN(_09022_));
 AND2_X1 _18679_ (.A1(_09020_),
    .A2(_08852_),
    .ZN(_09023_));
 NOR2_X1 _18680_ (.A1(_09022_),
    .A2(_09023_),
    .ZN(_09024_));
 AND2_X1 _18681_ (.A1(_08864_),
    .A2(_09002_),
    .ZN(_09025_));
 CLKBUF_X2 _18682_ (.A(_09025_),
    .Z(_09026_));
 AND2_X1 _18683_ (.A1(_09026_),
    .A2(_08965_),
    .ZN(_09027_));
 INV_X1 _18684_ (.A(_09027_),
    .ZN(_09028_));
 BUF_X2 _18685_ (.A(_08874_),
    .Z(_09029_));
 OAI221_X1 _18686_ (.A(_09026_),
    .B1(_08844_),
    .B2(_08845_),
    .C1(_09029_),
    .C2(_08843_),
    .ZN(_09030_));
 BUF_X2 _18687_ (.A(_09020_),
    .Z(_09031_));
 OAI21_X1 _18688_ (.A(_09031_),
    .B1(_08821_),
    .B2(_08989_),
    .ZN(_09032_));
 AND4_X1 _18689_ (.A1(_09024_),
    .A2(_09028_),
    .A3(_09030_),
    .A4(_09032_),
    .ZN(_09033_));
 NAND4_X2 _18690_ (.A1(_08975_),
    .A2(_09001_),
    .A3(_09019_),
    .A4(_09033_),
    .ZN(_09034_));
 NOR2_X4 _18691_ (.A1(_08948_),
    .A2(_09034_),
    .ZN(_09035_));
 XNOR2_X1 _18692_ (.A(_08815_),
    .B(_09035_),
    .ZN(_09036_));
 XNOR2_X1 _18693_ (.A(_09036_),
    .B(_04132_),
    .ZN(_09037_));
 INV_X2 _18694_ (.A(_01331_),
    .ZN(_09038_));
 BUF_X2 _18695_ (.A(_09038_),
    .Z(_09039_));
 BUF_X2 _18696_ (.A(_09039_),
    .Z(_09040_));
 MUX2_X1 _18697_ (.A(_04143_),
    .B(_09037_),
    .S(_09040_),
    .Z(_00724_));
 BUF_X2 _18698_ (.A(_17078_),
    .Z(_09041_));
 XOR2_X1 _18699_ (.A(_09041_),
    .B(_16974_),
    .Z(_09042_));
 AND2_X1 _18700_ (.A1(_08976_),
    .A2(_08902_),
    .ZN(_09043_));
 AND2_X1 _18701_ (.A1(_08976_),
    .A2(_08968_),
    .ZN(_09044_));
 OR2_X1 _18702_ (.A1(_09043_),
    .A2(_09044_),
    .ZN(_09045_));
 AND2_X1 _18703_ (.A1(_08849_),
    .A2(_08964_),
    .ZN(_09046_));
 AOI221_X1 _18704_ (.A(_09045_),
    .B1(_09046_),
    .B2(_08976_),
    .C1(_08821_),
    .C2(_09020_),
    .ZN(_09047_));
 AND2_X1 _18705_ (.A1(_08835_),
    .A2(_08822_),
    .ZN(_09048_));
 NAND3_X1 _18706_ (.A1(_08900_),
    .A2(_08845_),
    .A3(_09048_),
    .ZN(_09049_));
 AND2_X2 _18707_ (.A1(_08817_),
    .A2(_08964_),
    .ZN(_09050_));
 NAND2_X1 _18708_ (.A1(_09025_),
    .A2(_09050_),
    .ZN(_09051_));
 NAND2_X1 _18709_ (.A1(_09049_),
    .A2(_09051_),
    .ZN(_09052_));
 CLKBUF_X2 _18710_ (.A(_08957_),
    .Z(_09053_));
 AOI221_X4 _18711_ (.A(_09052_),
    .B1(_09020_),
    .B2(_09009_),
    .C1(_09053_),
    .C2(_08838_),
    .ZN(_09054_));
 AND4_X1 _18712_ (.A1(_08876_),
    .A2(_09047_),
    .A3(_08871_),
    .A4(_09054_),
    .ZN(_09055_));
 INV_X1 _18713_ (.A(_09050_),
    .ZN(_09056_));
 INV_X1 _18714_ (.A(_08834_),
    .ZN(_09057_));
 OAI221_X1 _18715_ (.A(_08953_),
    .B1(_09056_),
    .B2(_08995_),
    .C1(_09057_),
    .C2(_08991_),
    .ZN(_09058_));
 AND2_X1 _18716_ (.A1(_08987_),
    .A2(_08829_),
    .ZN(_09059_));
 AND2_X1 _18717_ (.A1(_08853_),
    .A2(_08828_),
    .ZN(_09060_));
 NAND2_X1 _18718_ (.A1(_08867_),
    .A2(_08877_),
    .ZN(_09061_));
 INV_X1 _18719_ (.A(_09061_),
    .ZN(_09062_));
 AND3_X1 _18720_ (.A1(_09062_),
    .A2(_08847_),
    .A3(_08873_),
    .ZN(_09063_));
 NOR4_X1 _18721_ (.A1(_09058_),
    .A2(_09059_),
    .A3(_09060_),
    .A4(_09063_),
    .ZN(_09064_));
 NAND3_X1 _18722_ (.A1(_08919_),
    .A2(_08867_),
    .A3(_08830_),
    .ZN(_09065_));
 NAND2_X1 _18723_ (.A1(_08830_),
    .A2(_08915_),
    .ZN(_09066_));
 NAND2_X1 _18724_ (.A1(_08986_),
    .A2(_08830_),
    .ZN(_09067_));
 AND4_X1 _18725_ (.A1(_08922_),
    .A2(_09065_),
    .A3(_09066_),
    .A4(_09067_),
    .ZN(_09068_));
 AND2_X1 _18726_ (.A1(_08834_),
    .A2(_09046_),
    .ZN(_09069_));
 AND2_X1 _18727_ (.A1(_08834_),
    .A2(_08969_),
    .ZN(_09070_));
 NOR2_X1 _18728_ (.A1(_09069_),
    .A2(_09070_),
    .ZN(_09071_));
 AND2_X1 _18729_ (.A1(_08887_),
    .A2(_08855_),
    .ZN(_09072_));
 AND2_X1 _18730_ (.A1(_08865_),
    .A2(_08908_),
    .ZN(_09073_));
 NOR2_X1 _18731_ (.A1(_09061_),
    .A2(_08964_),
    .ZN(_09074_));
 BUF_X2 _18732_ (.A(_08865_),
    .Z(_09075_));
 AOI211_X1 _18733_ (.A(_09072_),
    .B(_09073_),
    .C1(_09074_),
    .C2(_09075_),
    .ZN(_09076_));
 AND2_X2 _18734_ (.A1(_08877_),
    .A2(_16791_),
    .ZN(_09077_));
 AOI22_X1 _18735_ (.A1(_09077_),
    .A2(_08901_),
    .B1(_08929_),
    .B2(_08987_),
    .ZN(_09078_));
 AOI22_X1 _18736_ (.A1(_08941_),
    .A2(_08989_),
    .B1(_09008_),
    .B2(_08909_),
    .ZN(_09079_));
 AND4_X1 _18737_ (.A1(_09071_),
    .A2(_09076_),
    .A3(_09078_),
    .A4(_09079_),
    .ZN(_09080_));
 NAND4_X1 _18738_ (.A1(_09055_),
    .A2(_09064_),
    .A3(_09068_),
    .A4(_09080_),
    .ZN(_09081_));
 OAI21_X1 _18739_ (.A(_08941_),
    .B1(_09021_),
    .B2(_08855_),
    .ZN(_09082_));
 NAND4_X1 _18740_ (.A1(_08914_),
    .A2(_08973_),
    .A3(_09029_),
    .A4(_08827_),
    .ZN(_09083_));
 NAND2_X1 _18741_ (.A1(_09082_),
    .A2(_09083_),
    .ZN(_09084_));
 OAI21_X1 _18742_ (.A(_08982_),
    .B1(_09017_),
    .B2(_08945_),
    .ZN(_09085_));
 OAI21_X1 _18743_ (.A(_09085_),
    .B1(_08999_),
    .B2(_08983_),
    .ZN(_09086_));
 BUF_X2 _18744_ (.A(_08994_),
    .Z(_09087_));
 NOR2_X1 _18745_ (.A1(_08845_),
    .A2(_16793_),
    .ZN(_09088_));
 AOI211_X1 _18746_ (.A(_09084_),
    .B(_09086_),
    .C1(_09087_),
    .C2(_09088_),
    .ZN(_09089_));
 OAI21_X1 _18747_ (.A(_09026_),
    .B1(_08860_),
    .B2(_08855_),
    .ZN(_09090_));
 NAND3_X1 _18748_ (.A1(_08907_),
    .A2(_09003_),
    .A3(_08913_),
    .ZN(_09091_));
 AND2_X1 _18749_ (.A1(_09090_),
    .A2(_09091_),
    .ZN(_09092_));
 AND2_X2 _18750_ (.A1(_08874_),
    .A2(_16791_),
    .ZN(_09093_));
 OAI21_X1 _18751_ (.A(_09005_),
    .B1(_09093_),
    .B2(_09048_),
    .ZN(_09094_));
 NOR2_X2 _18752_ (.A1(_08918_),
    .A2(_08858_),
    .ZN(_09095_));
 OAI21_X1 _18753_ (.A(_08972_),
    .B1(_09095_),
    .B2(_08986_),
    .ZN(_09096_));
 INV_X1 _18754_ (.A(_09031_),
    .ZN(_09097_));
 NAND2_X1 _18755_ (.A1(_08824_),
    .A2(_08868_),
    .ZN(_09098_));
 NOR2_X1 _18756_ (.A1(_09097_),
    .A2(_09098_),
    .ZN(_09099_));
 INV_X1 _18757_ (.A(_09099_),
    .ZN(_09100_));
 NAND4_X1 _18758_ (.A1(_09092_),
    .A2(_09094_),
    .A3(_09096_),
    .A4(_09100_),
    .ZN(_09101_));
 AND3_X1 _18759_ (.A1(_08919_),
    .A2(_08900_),
    .A3(_08867_),
    .ZN(_09102_));
 AND2_X1 _18760_ (.A1(_08821_),
    .A2(_09004_),
    .ZN(_09103_));
 AND3_X1 _18761_ (.A1(_08968_),
    .A2(_08886_),
    .A3(_08899_),
    .ZN(_09104_));
 OR3_X1 _18762_ (.A1(_09102_),
    .A2(_09103_),
    .A3(_09104_),
    .ZN(_09105_));
 BUF_X2 _18763_ (.A(_08906_),
    .Z(_09106_));
 CLKBUF_X2 _18764_ (.A(_08877_),
    .Z(_09107_));
 OAI21_X1 _18765_ (.A(_09106_),
    .B1(_08889_),
    .B2(_09107_),
    .ZN(_09108_));
 INV_X1 _18766_ (.A(_09004_),
    .ZN(_09109_));
 OAI21_X1 _18767_ (.A(_09108_),
    .B1(_09109_),
    .B2(_08918_),
    .ZN(_09110_));
 NAND2_X1 _18768_ (.A1(_08873_),
    .A2(_08868_),
    .ZN(_09111_));
 NOR2_X1 _18769_ (.A1(_08892_),
    .A2(_09111_),
    .ZN(_09112_));
 INV_X1 _18770_ (.A(_09112_),
    .ZN(_09113_));
 OAI21_X1 _18771_ (.A(_08929_),
    .B1(_09093_),
    .B2(_08860_),
    .ZN(_09114_));
 CLKBUF_X2 _18772_ (.A(_08820_),
    .Z(_09115_));
 INV_X1 _18773_ (.A(_09115_),
    .ZN(_09116_));
 NAND3_X1 _18774_ (.A1(_08929_),
    .A2(_08868_),
    .A3(_09116_),
    .ZN(_09117_));
 NOR3_X1 _18775_ (.A1(_09115_),
    .A2(_08848_),
    .A3(_16793_),
    .ZN(_09118_));
 NAND3_X1 _18776_ (.A1(_09118_),
    .A2(_08913_),
    .A3(_08914_),
    .ZN(_09119_));
 NAND4_X1 _18777_ (.A1(_09113_),
    .A2(_09114_),
    .A3(_09117_),
    .A4(_09119_),
    .ZN(_09120_));
 NOR4_X1 _18778_ (.A1(_09101_),
    .A2(_09105_),
    .A3(_09110_),
    .A4(_09120_),
    .ZN(_09121_));
 INV_X1 _18779_ (.A(_09111_),
    .ZN(_09122_));
 NAND3_X1 _18780_ (.A1(_09122_),
    .A2(_08867_),
    .A3(_09008_),
    .ZN(_09123_));
 AND2_X1 _18781_ (.A1(_08855_),
    .A2(_08957_),
    .ZN(_09124_));
 AOI221_X4 _18782_ (.A(_09124_),
    .B1(_08852_),
    .B2(_08951_),
    .C1(_09053_),
    .C2(_09093_),
    .ZN(_09125_));
 AND2_X1 _18783_ (.A1(_08904_),
    .A2(_08952_),
    .ZN(_09126_));
 INV_X1 _18784_ (.A(_09126_),
    .ZN(_09127_));
 OAI21_X1 _18785_ (.A(_08848_),
    .B1(_08873_),
    .B2(_16793_),
    .ZN(_09128_));
 AND3_X1 _18786_ (.A1(_08825_),
    .A2(_08827_),
    .A3(_08848_),
    .ZN(_09129_));
 AOI22_X1 _18787_ (.A1(_09128_),
    .A2(_09129_),
    .B1(_08904_),
    .B2(_08994_),
    .ZN(_09130_));
 AND4_X1 _18788_ (.A1(_09123_),
    .A2(_09125_),
    .A3(_09127_),
    .A4(_09130_),
    .ZN(_09131_));
 AOI22_X1 _18789_ (.A1(_08887_),
    .A2(_08954_),
    .B1(_08907_),
    .B2(_08829_),
    .ZN(_09132_));
 NAND2_X1 _18790_ (.A1(_08865_),
    .A2(_09009_),
    .ZN(_09133_));
 OAI211_X1 _18791_ (.A(_09132_),
    .B(_09133_),
    .C1(_09057_),
    .C2(_09015_),
    .ZN(_09134_));
 NAND2_X1 _18792_ (.A1(_09106_),
    .A2(_09021_),
    .ZN(_09135_));
 NAND2_X1 _18793_ (.A1(_08940_),
    .A2(_09050_),
    .ZN(_09136_));
 NAND2_X1 _18794_ (.A1(_09046_),
    .A2(_08887_),
    .ZN(_09137_));
 NAND2_X1 _18795_ (.A1(_08860_),
    .A2(_08887_),
    .ZN(_09138_));
 NAND4_X1 _18796_ (.A1(_09135_),
    .A2(_09136_),
    .A3(_09137_),
    .A4(_09138_),
    .ZN(_09139_));
 AND2_X1 _18797_ (.A1(_08943_),
    .A2(_08994_),
    .ZN(_09140_));
 NAND2_X1 _18798_ (.A1(_09021_),
    .A2(_08994_),
    .ZN(_09141_));
 INV_X1 _18799_ (.A(_09021_),
    .ZN(_09142_));
 INV_X1 _18800_ (.A(_08957_),
    .ZN(_09143_));
 OAI21_X1 _18801_ (.A(_09141_),
    .B1(_09142_),
    .B2(_09143_),
    .ZN(_09144_));
 NOR4_X1 _18802_ (.A1(_09134_),
    .A2(_09139_),
    .A3(_09140_),
    .A4(_09144_),
    .ZN(_09145_));
 NAND4_X1 _18803_ (.A1(_09089_),
    .A2(_09121_),
    .A3(_09131_),
    .A4(_09145_),
    .ZN(_09146_));
 NOR2_X2 _18804_ (.A1(_09081_),
    .A2(_09146_),
    .ZN(_09147_));
 XOR2_X2 _18805_ (.A(_09147_),
    .B(_09035_),
    .Z(_09148_));
 AND2_X1 _18806_ (.A1(_05118_),
    .A2(_04384_),
    .ZN(_09149_));
 AND2_X1 _18807_ (.A1(_09149_),
    .A2(_05401_),
    .ZN(_09150_));
 AND2_X1 _18808_ (.A1(_04395_),
    .A2(_05390_),
    .ZN(_09151_));
 AND4_X1 _18809_ (.A1(_04680_),
    .A2(_04658_),
    .A3(_05110_),
    .A4(_04833_),
    .ZN(_09152_));
 OR3_X1 _18810_ (.A1(_09150_),
    .A2(_09151_),
    .A3(_09152_),
    .ZN(_09153_));
 NAND4_X1 _18811_ (.A1(_05324_),
    .A2(_05192_),
    .A3(_04833_),
    .A4(_04950_),
    .ZN(_09154_));
 INV_X1 _18812_ (.A(_04263_),
    .ZN(_09155_));
 OAI21_X1 _18813_ (.A(_09154_),
    .B1(_09155_),
    .B2(_05423_),
    .ZN(_09156_));
 OR2_X1 _18814_ (.A1(_09153_),
    .A2(_09156_),
    .ZN(_09157_));
 BUF_X2 _18815_ (.A(_05687_),
    .Z(_09158_));
 AND3_X1 _18816_ (.A1(_05676_),
    .A2(_09158_),
    .A3(_05324_),
    .ZN(_09159_));
 AND2_X1 _18817_ (.A1(_05214_),
    .A2(_05797_),
    .ZN(_09160_));
 AND2_X1 _18818_ (.A1(_05214_),
    .A2(_04537_),
    .ZN(_09161_));
 AND2_X1 _18819_ (.A1(_05214_),
    .A2(_04307_),
    .ZN(_09162_));
 OR4_X1 _18820_ (.A1(_09159_),
    .A2(_09160_),
    .A3(_09161_),
    .A4(_09162_),
    .ZN(_09163_));
 NAND2_X1 _18821_ (.A1(_05379_),
    .A2(_05511_),
    .ZN(_09164_));
 NAND4_X1 _18822_ (.A1(_05368_),
    .A2(_05324_),
    .A3(_04439_),
    .A4(_04592_),
    .ZN(_09165_));
 AND2_X1 _18823_ (.A1(_09164_),
    .A2(_09165_),
    .ZN(_09166_));
 NAND2_X1 _18824_ (.A1(_05511_),
    .A2(_05092_),
    .ZN(_09167_));
 INV_X1 _18825_ (.A(_05522_),
    .ZN(_09168_));
 AND2_X1 _18826_ (.A1(_06468_),
    .A2(_04899_),
    .ZN(_09169_));
 INV_X1 _18827_ (.A(_09169_),
    .ZN(_09170_));
 OAI211_X1 _18828_ (.A(_09166_),
    .B(_09167_),
    .C1(_09168_),
    .C2(_09170_),
    .ZN(_09171_));
 AND2_X1 _18829_ (.A1(_04537_),
    .A2(_05291_),
    .ZN(_09172_));
 AND2_X1 _18830_ (.A1(_05291_),
    .A2(_04559_),
    .ZN(_09173_));
 NOR2_X1 _18831_ (.A1(_09172_),
    .A2(_09173_),
    .ZN(_09174_));
 AND2_X1 _18832_ (.A1(_05258_),
    .A2(_05120_),
    .ZN(_09175_));
 INV_X1 _18833_ (.A(_09175_),
    .ZN(_09176_));
 NAND2_X1 _18834_ (.A1(_05291_),
    .A2(_05225_),
    .ZN(_09177_));
 BUF_X2 _18835_ (.A(_05709_),
    .Z(_09178_));
 NAND2_X1 _18836_ (.A1(_09178_),
    .A2(_05291_),
    .ZN(_09179_));
 NAND4_X1 _18837_ (.A1(_09174_),
    .A2(_09176_),
    .A3(_09177_),
    .A4(_09179_),
    .ZN(_09180_));
 NOR4_X1 _18838_ (.A1(_09157_),
    .A2(_09163_),
    .A3(_09171_),
    .A4(_09180_),
    .ZN(_09181_));
 AND2_X2 _18839_ (.A1(_04658_),
    .A2(_05137_),
    .ZN(_09182_));
 INV_X1 _18840_ (.A(_09182_),
    .ZN(_09183_));
 AOI21_X1 _18841_ (.A(_04800_),
    .B1(_04526_),
    .B2(_09183_),
    .ZN(_09184_));
 INV_X1 _18842_ (.A(_09149_),
    .ZN(_09185_));
 INV_X1 _18843_ (.A(_04395_),
    .ZN(_09186_));
 AOI21_X1 _18844_ (.A(_04800_),
    .B1(_09185_),
    .B2(_09186_),
    .ZN(_09187_));
 NAND2_X1 _18845_ (.A1(_06226_),
    .A2(_04614_),
    .ZN(_09188_));
 INV_X1 _18846_ (.A(_04450_),
    .ZN(_09189_));
 OAI21_X1 _18847_ (.A(_09188_),
    .B1(_09189_),
    .B2(_04800_),
    .ZN(_09190_));
 NOR3_X1 _18848_ (.A1(_09184_),
    .A2(_09187_),
    .A3(_09190_),
    .ZN(_09191_));
 AND2_X1 _18849_ (.A1(_04844_),
    .A2(_04921_),
    .ZN(_09192_));
 INV_X1 _18850_ (.A(_04844_),
    .ZN(_09193_));
 INV_X1 _18851_ (.A(_04746_),
    .ZN(_09194_));
 AOI21_X1 _18852_ (.A(_09193_),
    .B1(_09189_),
    .B2(_09194_),
    .ZN(_09195_));
 AOI211_X1 _18853_ (.A(_09192_),
    .B(_09195_),
    .C1(_04888_),
    .C2(_09169_),
    .ZN(_09196_));
 INV_X2 _18854_ (.A(_04997_),
    .ZN(_09197_));
 INV_X1 _18855_ (.A(_04340_),
    .ZN(_09198_));
 AOI21_X1 _18856_ (.A(_09197_),
    .B1(_09198_),
    .B2(_05456_),
    .ZN(_09199_));
 INV_X1 _18857_ (.A(_05478_),
    .ZN(_09200_));
 INV_X1 _18858_ (.A(_05096_),
    .ZN(_09201_));
 AOI21_X1 _18859_ (.A(_09197_),
    .B1(_09200_),
    .B2(_09201_),
    .ZN(_09202_));
 AND2_X1 _18860_ (.A1(_05045_),
    .A2(_04537_),
    .ZN(_09203_));
 AND2_X1 _18861_ (.A1(_05045_),
    .A2(_05599_),
    .ZN(_09204_));
 NOR4_X1 _18862_ (.A1(_09199_),
    .A2(_09202_),
    .A3(_09203_),
    .A4(_09204_),
    .ZN(_09205_));
 AND2_X1 _18863_ (.A1(_06534_),
    .A2(_04494_),
    .ZN(_09206_));
 AND4_X1 _18864_ (.A1(_05192_),
    .A2(_04461_),
    .A3(_04713_),
    .A4(_04472_),
    .ZN(_09207_));
 AND4_X1 _18865_ (.A1(_05137_),
    .A2(_04461_),
    .A3(_04669_),
    .A4(_04472_),
    .ZN(_09208_));
 NOR4_X1 _18866_ (.A1(_09206_),
    .A2(_04406_),
    .A3(_09207_),
    .A4(_09208_),
    .ZN(_09209_));
 AND4_X1 _18867_ (.A1(_09191_),
    .A2(_09196_),
    .A3(_09205_),
    .A4(_09209_),
    .ZN(_09210_));
 AND3_X1 _18868_ (.A1(_06281_),
    .A2(_06303_),
    .A3(_05313_),
    .ZN(_09211_));
 AND3_X1 _18869_ (.A1(_06270_),
    .A2(_04713_),
    .A3(_04735_),
    .ZN(_09212_));
 AND3_X1 _18870_ (.A1(_06270_),
    .A2(_04713_),
    .A3(_05368_),
    .ZN(_09213_));
 NOR3_X1 _18871_ (.A1(_09211_),
    .A2(_09212_),
    .A3(_09213_),
    .ZN(_09214_));
 AND2_X1 _18872_ (.A1(_04559_),
    .A2(_06281_),
    .ZN(_09215_));
 AND3_X1 _18873_ (.A1(_06270_),
    .A2(_05368_),
    .A3(_04658_),
    .ZN(_09216_));
 NOR2_X1 _18874_ (.A1(_09215_),
    .A2(_09216_),
    .ZN(_09217_));
 OAI21_X1 _18875_ (.A(_06281_),
    .B1(_04636_),
    .B2(_05159_),
    .ZN(_09218_));
 NAND4_X1 _18876_ (.A1(_09214_),
    .A2(_06358_),
    .A3(_09217_),
    .A4(_09218_),
    .ZN(_09219_));
 AND2_X1 _18877_ (.A1(_06226_),
    .A2(_06391_),
    .ZN(_09220_));
 INV_X1 _18878_ (.A(_09220_),
    .ZN(_09221_));
 OAI211_X1 _18879_ (.A(_06446_),
    .B(_04950_),
    .C1(_06314_),
    .C2(_05203_),
    .ZN(_09222_));
 NAND2_X1 _18880_ (.A1(_09221_),
    .A2(_09222_),
    .ZN(_09223_));
 AND2_X1 _18881_ (.A1(_06160_),
    .A2(_09182_),
    .ZN(_09224_));
 INV_X1 _18882_ (.A(_09224_),
    .ZN(_09225_));
 AND2_X1 _18883_ (.A1(_06171_),
    .A2(_04395_),
    .ZN(_09226_));
 INV_X1 _18884_ (.A(_09226_),
    .ZN(_09227_));
 AND2_X1 _18885_ (.A1(_04713_),
    .A2(_05116_),
    .ZN(_09228_));
 OAI21_X1 _18886_ (.A(_06171_),
    .B1(_09228_),
    .B2(_04778_),
    .ZN(_09229_));
 NAND3_X1 _18887_ (.A1(_09225_),
    .A2(_09227_),
    .A3(_09229_),
    .ZN(_09230_));
 OAI211_X1 _18888_ (.A(_06567_),
    .B(_05863_),
    .C1(_04959_),
    .C2(_06325_),
    .ZN(_09231_));
 OAI211_X1 _18889_ (.A(_06567_),
    .B(_05797_),
    .C1(_04959_),
    .C2(_05192_),
    .ZN(_09232_));
 NAND3_X1 _18890_ (.A1(_06567_),
    .A2(_06325_),
    .A3(_06303_),
    .ZN(_09233_));
 NAND4_X1 _18891_ (.A1(_06578_),
    .A2(_09231_),
    .A3(_09232_),
    .A4(_09233_),
    .ZN(_09234_));
 NOR4_X1 _18892_ (.A1(_09219_),
    .A2(_09223_),
    .A3(_09230_),
    .A4(_09234_),
    .ZN(_09235_));
 OAI21_X1 _18893_ (.A(_05786_),
    .B1(_05929_),
    .B2(_04855_),
    .ZN(_09236_));
 OAI211_X1 _18894_ (.A(_05786_),
    .B(_05797_),
    .C1(_06314_),
    .C2(_05203_),
    .ZN(_09237_));
 INV_X2 _18895_ (.A(_05775_),
    .ZN(_09238_));
 OAI211_X1 _18896_ (.A(_09236_),
    .B(_09237_),
    .C1(_06105_),
    .C2(_09238_),
    .ZN(_09239_));
 NAND4_X1 _18897_ (.A1(_09158_),
    .A2(_06325_),
    .A3(_05874_),
    .A4(_04950_),
    .ZN(_09240_));
 OAI21_X1 _18898_ (.A(_05632_),
    .B1(_09178_),
    .B2(_05064_),
    .ZN(_09241_));
 OAI211_X1 _18899_ (.A(_09158_),
    .B(_05874_),
    .C1(_05096_),
    .C2(_06490_),
    .ZN(_09242_));
 NAND4_X1 _18900_ (.A1(_05621_),
    .A2(_09240_),
    .A3(_09241_),
    .A4(_09242_),
    .ZN(_09243_));
 AND2_X1 _18901_ (.A1(_04296_),
    .A2(_06017_),
    .ZN(_09244_));
 INV_X1 _18902_ (.A(_09244_),
    .ZN(_09245_));
 BUF_X2 _18903_ (.A(_06017_),
    .Z(_09246_));
 OAI21_X1 _18904_ (.A(_09246_),
    .B1(_04559_),
    .B2(_05159_),
    .ZN(_09247_));
 INV_X1 _18905_ (.A(_06017_),
    .ZN(_09248_));
 OAI211_X1 _18906_ (.A(_09245_),
    .B(_09247_),
    .C1(_09155_),
    .C2(_09248_),
    .ZN(_09249_));
 OAI211_X1 _18907_ (.A(_05907_),
    .B(_05863_),
    .C1(_04959_),
    .C2(_05192_),
    .ZN(_09250_));
 BUF_X2 _18908_ (.A(_05896_),
    .Z(_09251_));
 NAND2_X1 _18909_ (.A1(_04263_),
    .A2(_09251_),
    .ZN(_09252_));
 NAND3_X1 _18910_ (.A1(_05096_),
    .A2(_04472_),
    .A3(_05874_),
    .ZN(_09253_));
 NAND3_X1 _18911_ (.A1(_09251_),
    .A2(_05203_),
    .A3(_04636_),
    .ZN(_09254_));
 NAND4_X1 _18912_ (.A1(_09250_),
    .A2(_09252_),
    .A3(_09253_),
    .A4(_09254_),
    .ZN(_09255_));
 NOR4_X1 _18913_ (.A1(_09239_),
    .A2(_09243_),
    .A3(_09249_),
    .A4(_09255_),
    .ZN(_09256_));
 NAND4_X1 _18914_ (.A1(_09181_),
    .A2(_09210_),
    .A3(_09235_),
    .A4(_09256_),
    .ZN(_09257_));
 NOR2_X2 _18915_ (.A1(_09257_),
    .A2(_06672_),
    .ZN(_09258_));
 XNOR2_X1 _18916_ (.A(_09148_),
    .B(_09258_),
    .ZN(_09259_));
 AND2_X1 _18917_ (.A1(_06941_),
    .A2(_07565_),
    .ZN(_09260_));
 INV_X2 _18918_ (.A(_07565_),
    .ZN(_09261_));
 AND2_X1 _18919_ (.A1(_16712_),
    .A2(_16714_),
    .ZN(_09262_));
 AND2_X1 _18920_ (.A1(_09262_),
    .A2(_16713_),
    .ZN(_09263_));
 INV_X1 _18921_ (.A(_09263_),
    .ZN(_09264_));
 AOI21_X1 _18922_ (.A(_09261_),
    .B1(_07959_),
    .B2(_09264_),
    .ZN(_09265_));
 AOI211_X1 _18923_ (.A(_09260_),
    .B(_09265_),
    .C1(_07795_),
    .C2(_07576_),
    .ZN(_09266_));
 OAI211_X1 _18924_ (.A(_08450_),
    .B(_08461_),
    .C1(_08459_),
    .C2(_07161_),
    .ZN(_09267_));
 OAI21_X1 _18925_ (.A(_06996_),
    .B1(_07609_),
    .B2(_07348_),
    .ZN(_09268_));
 NAND2_X1 _18926_ (.A1(_07795_),
    .A2(_08450_),
    .ZN(_09269_));
 NAND4_X1 _18927_ (.A1(_09266_),
    .A2(_09267_),
    .A3(_09268_),
    .A4(_09269_),
    .ZN(_09270_));
 OAI21_X1 _18928_ (.A(_08491_),
    .B1(_08308_),
    .B2(_08167_),
    .ZN(_09271_));
 AND2_X1 _18929_ (.A1(_06743_),
    .A2(_08091_),
    .ZN(_09272_));
 INV_X1 _18930_ (.A(_09272_),
    .ZN(_09273_));
 OAI21_X1 _18931_ (.A(_09271_),
    .B1(_08492_),
    .B2(_09273_),
    .ZN(_09274_));
 NAND3_X1 _18932_ (.A1(_07348_),
    .A2(_08189_),
    .A3(_07543_),
    .ZN(_09275_));
 NAND4_X1 _18933_ (.A1(_08200_),
    .A2(_07150_),
    .A3(_08461_),
    .A4(_07543_),
    .ZN(_09276_));
 INV_X1 _18934_ (.A(_07609_),
    .ZN(_09277_));
 OAI211_X1 _18935_ (.A(_09275_),
    .B(_09276_),
    .C1(_08492_),
    .C2(_09277_),
    .ZN(_09278_));
 OAI21_X1 _18936_ (.A(_07249_),
    .B1(_08454_),
    .B2(_08498_),
    .ZN(_09279_));
 AND2_X1 _18937_ (.A1(_07948_),
    .A2(_07238_),
    .ZN(_09280_));
 INV_X1 _18938_ (.A(_09280_),
    .ZN(_09281_));
 AND2_X1 _18939_ (.A1(_07337_),
    .A2(_07238_),
    .ZN(_09282_));
 INV_X1 _18940_ (.A(_09282_),
    .ZN(_09283_));
 NAND2_X1 _18941_ (.A1(_07227_),
    .A2(_09263_),
    .ZN(_09284_));
 NAND4_X1 _18942_ (.A1(_09279_),
    .A2(_09281_),
    .A3(_09283_),
    .A4(_09284_),
    .ZN(_09285_));
 NOR4_X1 _18943_ (.A1(_09270_),
    .A2(_09274_),
    .A3(_09278_),
    .A4(_09285_),
    .ZN(_09286_));
 NAND2_X2 _18944_ (.A1(_09262_),
    .A2(_06908_),
    .ZN(_09287_));
 INV_X1 _18945_ (.A(_09287_),
    .ZN(_09288_));
 BUF_X2 _18946_ (.A(_09288_),
    .Z(_09289_));
 OAI21_X1 _18947_ (.A(_08025_),
    .B1(_08047_),
    .B2(_09289_),
    .ZN(_09290_));
 NAND4_X1 _18948_ (.A1(_08200_),
    .A2(_07194_),
    .A3(_07161_),
    .A4(_08463_),
    .ZN(_09291_));
 INV_X1 _18949_ (.A(_08014_),
    .ZN(_09292_));
 OAI211_X1 _18950_ (.A(_09290_),
    .B(_09291_),
    .C1(_07707_),
    .C2(_09292_),
    .ZN(_09293_));
 INV_X1 _18951_ (.A(_06787_),
    .ZN(_09294_));
 NAND2_X1 _18952_ (.A1(_07378_),
    .A2(_06732_),
    .ZN(_09295_));
 AND2_X1 _18953_ (.A1(_08431_),
    .A2(_07183_),
    .ZN(_09296_));
 NAND2_X1 _18954_ (.A1(_09296_),
    .A2(_06732_),
    .ZN(_09297_));
 NAND2_X1 _18955_ (.A1(_06732_),
    .A2(_09262_),
    .ZN(_09298_));
 NAND4_X1 _18956_ (.A1(_09294_),
    .A2(_09295_),
    .A3(_09297_),
    .A4(_09298_),
    .ZN(_09299_));
 OAI211_X1 _18957_ (.A(_07411_),
    .B(_08461_),
    .C1(_08459_),
    .C2(_08102_),
    .ZN(_09300_));
 OAI211_X1 _18958_ (.A(_07411_),
    .B(_08233_),
    .C1(_08459_),
    .C2(_07161_),
    .ZN(_09301_));
 NAND2_X1 _18959_ (.A1(_08498_),
    .A2(_07411_),
    .ZN(_09302_));
 NAND4_X1 _18960_ (.A1(_09300_),
    .A2(_09301_),
    .A3(_08474_),
    .A4(_09302_),
    .ZN(_09303_));
 INV_X1 _18961_ (.A(_07828_),
    .ZN(_09304_));
 INV_X1 _18962_ (.A(_09296_),
    .ZN(_09305_));
 INV_X1 _18963_ (.A(_06886_),
    .ZN(_09306_));
 AOI21_X1 _18964_ (.A(_09304_),
    .B1(_09305_),
    .B2(_09306_),
    .ZN(_09307_));
 NOR4_X1 _18965_ (.A1(_09293_),
    .A2(_09299_),
    .A3(_09303_),
    .A4(_09307_),
    .ZN(_09308_));
 NAND2_X1 _18966_ (.A1(_07795_),
    .A2(_07893_),
    .ZN(_09309_));
 INV_X1 _18967_ (.A(_06941_),
    .ZN(_09310_));
 INV_X1 _18968_ (.A(_07893_),
    .ZN(_09311_));
 OAI21_X1 _18969_ (.A(_09309_),
    .B1(_09310_),
    .B2(_09311_),
    .ZN(_09312_));
 AND2_X2 _18970_ (.A1(_06864_),
    .A2(_07356_),
    .ZN(_09313_));
 INV_X1 _18971_ (.A(_09313_),
    .ZN(_09314_));
 AOI21_X1 _18972_ (.A(_09311_),
    .B1(_09314_),
    .B2(_08482_),
    .ZN(_09315_));
 NAND4_X1 _18973_ (.A1(_08069_),
    .A2(_08080_),
    .A3(_06930_),
    .A4(_06699_),
    .ZN(_09316_));
 OAI21_X1 _18974_ (.A(_09316_),
    .B1(_09287_),
    .B2(_09311_),
    .ZN(_09317_));
 AND4_X1 _18975_ (.A1(_08102_),
    .A2(_08080_),
    .A3(_08478_),
    .A4(_06699_),
    .ZN(_09318_));
 NOR4_X1 _18976_ (.A1(_09312_),
    .A2(_09315_),
    .A3(_09317_),
    .A4(_09318_),
    .ZN(_09319_));
 INV_X1 _18977_ (.A(_08156_),
    .ZN(_09320_));
 AND2_X2 _18978_ (.A1(_06919_),
    .A2(_07598_),
    .ZN(_09321_));
 INV_X1 _18979_ (.A(_09321_),
    .ZN(_09322_));
 AOI21_X1 _18980_ (.A(_09320_),
    .B1(_08453_),
    .B2(_09322_),
    .ZN(_09323_));
 NOR2_X1 _18981_ (.A1(_07740_),
    .A2(_07150_),
    .ZN(_09324_));
 INV_X1 _18982_ (.A(_06875_),
    .ZN(_09325_));
 AND3_X1 _18983_ (.A1(_08156_),
    .A2(_09324_),
    .A3(_09325_),
    .ZN(_09326_));
 AND2_X1 _18984_ (.A1(_07139_),
    .A2(_07117_),
    .ZN(_09327_));
 AND2_X1 _18985_ (.A1(_08145_),
    .A2(_09327_),
    .ZN(_09328_));
 NOR2_X1 _18986_ (.A1(_07106_),
    .A2(_16712_),
    .ZN(_09329_));
 AND2_X2 _18987_ (.A1(_09329_),
    .A2(_06908_),
    .ZN(_09330_));
 AND2_X1 _18988_ (.A1(_08145_),
    .A2(_09330_),
    .ZN(_09331_));
 NOR4_X1 _18989_ (.A1(_09323_),
    .A2(_09326_),
    .A3(_09328_),
    .A4(_09331_),
    .ZN(_09332_));
 OAI21_X1 _18990_ (.A(_07095_),
    .B1(_08047_),
    .B2(_09289_),
    .ZN(_09333_));
 NAND2_X1 _18991_ (.A1(_07095_),
    .A2(_08473_),
    .ZN(_09334_));
 NAND4_X1 _18992_ (.A1(_07194_),
    .A2(_06974_),
    .A3(_08080_),
    .A4(_07161_),
    .ZN(_09335_));
 AND3_X1 _18993_ (.A1(_09333_),
    .A2(_09334_),
    .A3(_09335_),
    .ZN(_09336_));
 AND3_X1 _18994_ (.A1(_07861_),
    .A2(_08431_),
    .A3(_08422_),
    .ZN(_09337_));
 AND2_X1 _18995_ (.A1(_08413_),
    .A2(_07674_),
    .ZN(_09338_));
 AND2_X1 _18996_ (.A1(_07674_),
    .A2(_09272_),
    .ZN(_09339_));
 AND4_X1 _18997_ (.A1(_07183_),
    .A2(_08080_),
    .A3(_08403_),
    .A4(_07554_),
    .ZN(_09340_));
 NOR4_X1 _18998_ (.A1(_09337_),
    .A2(_09338_),
    .A3(_09339_),
    .A4(_09340_),
    .ZN(_09341_));
 AND4_X1 _18999_ (.A1(_09319_),
    .A2(_09332_),
    .A3(_09336_),
    .A4(_09341_),
    .ZN(_09342_));
 NAND4_X1 _19000_ (.A1(_08222_),
    .A2(_08478_),
    .A3(_07150_),
    .A4(_08113_),
    .ZN(_09343_));
 AND2_X1 _19001_ (.A1(_07477_),
    .A2(_09343_),
    .ZN(_09344_));
 NAND2_X1 _19002_ (.A1(_07466_),
    .A2(_07609_),
    .ZN(_09345_));
 INV_X1 _19003_ (.A(_07466_),
    .ZN(_09346_));
 OAI21_X1 _19004_ (.A(_07117_),
    .B1(_06930_),
    .B2(_06853_),
    .ZN(_09347_));
 NOR2_X1 _19005_ (.A1(_09347_),
    .A2(_08403_),
    .ZN(_09348_));
 INV_X1 _19006_ (.A(_09348_),
    .ZN(_09349_));
 OAI211_X1 _19007_ (.A(_09344_),
    .B(_09345_),
    .C1(_09346_),
    .C2(_09349_),
    .ZN(_09350_));
 AND2_X1 _19008_ (.A1(_07992_),
    .A2(_06809_),
    .ZN(_09351_));
 CLKBUF_X2 _19009_ (.A(_09351_),
    .Z(_09352_));
 NAND2_X1 _19010_ (.A1(_09352_),
    .A2(_06952_),
    .ZN(_09353_));
 NAND3_X1 _19011_ (.A1(_07762_),
    .A2(_08200_),
    .A3(_08222_),
    .ZN(_09354_));
 NAND2_X1 _19012_ (.A1(_09353_),
    .A2(_09354_),
    .ZN(_09355_));
 AND2_X1 _19013_ (.A1(_09352_),
    .A2(_08233_),
    .ZN(_09356_));
 AND2_X1 _19014_ (.A1(_09352_),
    .A2(_09330_),
    .ZN(_09357_));
 OR3_X1 _19015_ (.A1(_09355_),
    .A2(_09356_),
    .A3(_09357_),
    .ZN(_09358_));
 NOR2_X1 _19016_ (.A1(_07128_),
    .A2(_07150_),
    .ZN(_09359_));
 AND2_X1 _19017_ (.A1(_09359_),
    .A2(_08485_),
    .ZN(_09360_));
 INV_X1 _19018_ (.A(_09360_),
    .ZN(_09361_));
 NAND2_X1 _19019_ (.A1(_07631_),
    .A2(_08308_),
    .ZN(_09362_));
 NAND2_X1 _19020_ (.A1(_08485_),
    .A2(_07532_),
    .ZN(_09363_));
 NAND2_X1 _19021_ (.A1(_08485_),
    .A2(_06776_),
    .ZN(_09364_));
 NAND4_X1 _19022_ (.A1(_09361_),
    .A2(_09362_),
    .A3(_09363_),
    .A4(_09364_),
    .ZN(_09365_));
 OAI21_X1 _19023_ (.A(_07315_),
    .B1(_09313_),
    .B2(_08047_),
    .ZN(_09366_));
 OAI21_X1 _19024_ (.A(_07315_),
    .B1(_07795_),
    .B2(_08479_),
    .ZN(_09367_));
 NAND4_X1 _19025_ (.A1(_08222_),
    .A2(_08102_),
    .A3(_08461_),
    .A4(_07554_),
    .ZN(_09368_));
 NAND3_X1 _19026_ (.A1(_09366_),
    .A2(_09367_),
    .A3(_09368_),
    .ZN(_09369_));
 NOR4_X1 _19027_ (.A1(_09350_),
    .A2(_09358_),
    .A3(_09365_),
    .A4(_09369_),
    .ZN(_09370_));
 NAND4_X1 _19028_ (.A1(_09286_),
    .A2(_09308_),
    .A3(_09342_),
    .A4(_09370_),
    .ZN(_09371_));
 NOR2_X2 _19029_ (.A1(_09371_),
    .A2(_07040_),
    .ZN(_09372_));
 INV_X1 _19030_ (.A(_08702_),
    .ZN(_09373_));
 AOI211_X1 _19031_ (.A(_08652_),
    .B(_09373_),
    .C1(_08590_),
    .C2(_08587_),
    .ZN(_09374_));
 NAND2_X1 _19032_ (.A1(_08704_),
    .A2(_08703_),
    .ZN(_09375_));
 NAND2_X1 _19033_ (.A1(_08702_),
    .A2(_08621_),
    .ZN(_09376_));
 INV_X1 _19034_ (.A(_08613_),
    .ZN(_09377_));
 OAI211_X1 _19035_ (.A(_09375_),
    .B(_09376_),
    .C1(_09373_),
    .C2(_09377_),
    .ZN(_09378_));
 AND4_X1 _19036_ (.A1(_08733_),
    .A2(_08618_),
    .A3(_08539_),
    .A4(_08675_),
    .ZN(_09379_));
 NOR3_X1 _19037_ (.A1(_09374_),
    .A2(_09378_),
    .A3(_09379_),
    .ZN(_09380_));
 AND4_X1 _19038_ (.A1(_08631_),
    .A2(_08509_),
    .A3(_08642_),
    .A4(_08675_),
    .ZN(_09381_));
 BUF_X2 _19039_ (.A(_16703_),
    .Z(_09382_));
 AOI211_X1 _19040_ (.A(_08669_),
    .B(_08524_),
    .C1(_09382_),
    .C2(_08794_),
    .ZN(_09383_));
 AOI211_X1 _19041_ (.A(_09381_),
    .B(_09383_),
    .C1(_08607_),
    .C2(_08646_),
    .ZN(_09384_));
 OAI211_X1 _19042_ (.A(_08513_),
    .B(_08637_),
    .C1(_08651_),
    .C2(_08794_),
    .ZN(_09385_));
 NAND3_X1 _19043_ (.A1(_08665_),
    .A2(_08592_),
    .A3(_08731_),
    .ZN(_09386_));
 NAND4_X1 _19044_ (.A1(_08615_),
    .A2(_09382_),
    .A3(_08675_),
    .A4(_08633_),
    .ZN(_09387_));
 AND4_X1 _19045_ (.A1(_08514_),
    .A2(_09385_),
    .A3(_09386_),
    .A4(_09387_),
    .ZN(_09388_));
 AND2_X1 _19046_ (.A1(_08676_),
    .A2(_08714_),
    .ZN(_09389_));
 INV_X1 _19047_ (.A(_08764_),
    .ZN(_09390_));
 AOI21_X1 _19048_ (.A(_08727_),
    .B1(_09390_),
    .B2(_08802_),
    .ZN(_09391_));
 AOI211_X1 _19049_ (.A(_09389_),
    .B(_09391_),
    .C1(_08677_),
    .C2(_08747_),
    .ZN(_09392_));
 AND4_X1 _19050_ (.A1(_09380_),
    .A2(_09384_),
    .A3(_09388_),
    .A4(_09392_),
    .ZN(_09393_));
 INV_X1 _19051_ (.A(_08602_),
    .ZN(_09394_));
 OAI211_X1 _19052_ (.A(_08622_),
    .B(_16706_),
    .C1(_08794_),
    .C2(_16705_),
    .ZN(_09395_));
 NAND3_X1 _19053_ (.A1(_08599_),
    .A2(_08574_),
    .A3(_08614_),
    .ZN(_09396_));
 NAND3_X1 _19054_ (.A1(_08598_),
    .A2(_08618_),
    .A3(_08614_),
    .ZN(_09397_));
 AND4_X1 _19055_ (.A1(_09394_),
    .A2(_09395_),
    .A3(_09396_),
    .A4(_09397_),
    .ZN(_09398_));
 AND2_X1 _19056_ (.A1(_08568_),
    .A2(_08541_),
    .ZN(_09399_));
 AND2_X1 _19057_ (.A1(_08517_),
    .A2(_08525_),
    .ZN(_09400_));
 INV_X1 _19058_ (.A(_09400_),
    .ZN(_09401_));
 OAI21_X1 _19059_ (.A(_08790_),
    .B1(_08793_),
    .B2(_09401_),
    .ZN(_09402_));
 AOI211_X1 _19060_ (.A(_09399_),
    .B(_09402_),
    .C1(_08708_),
    .C2(_08542_),
    .ZN(_09403_));
 AND2_X1 _19061_ (.A1(_08590_),
    .A2(_08517_),
    .ZN(_09404_));
 OAI21_X1 _19062_ (.A(_08586_),
    .B1(_09404_),
    .B2(_08611_),
    .ZN(_09405_));
 NAND2_X1 _19063_ (.A1(_08544_),
    .A2(_08636_),
    .ZN(_09406_));
 OAI211_X1 _19064_ (.A(_08625_),
    .B(_08631_),
    .C1(_08579_),
    .C2(_08574_),
    .ZN(_09407_));
 OAI211_X1 _19065_ (.A(_08625_),
    .B(_08637_),
    .C1(_08651_),
    .C2(_08574_),
    .ZN(_09408_));
 AND4_X1 _19066_ (.A1(_08628_),
    .A2(_09406_),
    .A3(_09407_),
    .A4(_09408_),
    .ZN(_09409_));
 AND4_X1 _19067_ (.A1(_09398_),
    .A2(_09403_),
    .A3(_09405_),
    .A4(_09409_),
    .ZN(_09410_));
 AOI21_X1 _19068_ (.A(_08560_),
    .B1(_08801_),
    .B2(_08802_),
    .ZN(_09411_));
 AOI21_X1 _19069_ (.A(_08560_),
    .B1(_08710_),
    .B2(_08694_),
    .ZN(_09412_));
 AND2_X1 _19070_ (.A1(_09404_),
    .A2(_08559_),
    .ZN(_09413_));
 AND4_X1 _19071_ (.A1(_08579_),
    .A2(_08632_),
    .A3(_08633_),
    .A4(_08593_),
    .ZN(_09414_));
 NOR4_X1 _19072_ (.A1(_09411_),
    .A2(_09412_),
    .A3(_09413_),
    .A4(_09414_),
    .ZN(_09415_));
 INV_X1 _19073_ (.A(_08663_),
    .ZN(_09416_));
 INV_X1 _19074_ (.A(_08758_),
    .ZN(_09417_));
 AOI21_X1 _19075_ (.A(_09416_),
    .B1(_09417_),
    .B2(_08680_),
    .ZN(_09418_));
 AOI21_X1 _19076_ (.A(_09416_),
    .B1(_09390_),
    .B2(_08802_),
    .ZN(_09419_));
 AOI211_X1 _19077_ (.A(_09418_),
    .B(_09419_),
    .C1(_08664_),
    .C2(_08747_),
    .ZN(_09420_));
 OAI21_X1 _19078_ (.A(_08551_),
    .B1(_16703_),
    .B2(_08507_),
    .ZN(_09421_));
 INV_X1 _19079_ (.A(_09421_),
    .ZN(_09422_));
 AND2_X1 _19080_ (.A1(_08564_),
    .A2(_09422_),
    .ZN(_09423_));
 OAI21_X1 _19081_ (.A(_08569_),
    .B1(_08767_),
    .B2(_08801_),
    .ZN(_09424_));
 AOI211_X1 _19082_ (.A(_09423_),
    .B(_09424_),
    .C1(_08565_),
    .C2(_09400_),
    .ZN(_09425_));
 AOI21_X1 _19083_ (.A(_08558_),
    .B1(_08520_),
    .B2(_09377_),
    .ZN(_09426_));
 AOI211_X1 _19084_ (.A(_08775_),
    .B(_09426_),
    .C1(_08549_),
    .C2(_08746_),
    .ZN(_09427_));
 AND4_X1 _19085_ (.A1(_09415_),
    .A2(_09420_),
    .A3(_09425_),
    .A4(_09427_),
    .ZN(_09428_));
 NAND2_X1 _19086_ (.A1(_08619_),
    .A2(_08572_),
    .ZN(_09429_));
 NAND4_X1 _19087_ (.A1(_08580_),
    .A2(_08512_),
    .A3(_08618_),
    .A4(_08593_),
    .ZN(_09430_));
 AND2_X1 _19088_ (.A1(_08687_),
    .A2(_09430_),
    .ZN(_09431_));
 OAI21_X1 _19089_ (.A(_08650_),
    .B1(_08746_),
    .B2(_08573_),
    .ZN(_09432_));
 OAI21_X1 _19090_ (.A(_08605_),
    .B1(_08594_),
    .B2(_08684_),
    .ZN(_09433_));
 OAI21_X1 _19091_ (.A(_08604_),
    .B1(_08578_),
    .B2(_08637_),
    .ZN(_09434_));
 AND4_X1 _19092_ (.A1(_09431_),
    .A2(_09432_),
    .A3(_09433_),
    .A4(_09434_),
    .ZN(_09435_));
 AND2_X1 _19093_ (.A1(_08571_),
    .A2(_08600_),
    .ZN(_09436_));
 AND2_X1 _19094_ (.A1(_08572_),
    .A2(_08688_),
    .ZN(_09437_));
 AOI211_X1 _19095_ (.A(_09436_),
    .B(_09437_),
    .C1(_08704_),
    .C2(_08572_),
    .ZN(_09438_));
 NAND4_X1 _19096_ (.A1(_08641_),
    .A2(_08579_),
    .A3(_08631_),
    .A4(_08642_),
    .ZN(_09439_));
 AND2_X1 _19097_ (.A1(_08608_),
    .A2(_08714_),
    .ZN(_09440_));
 INV_X1 _19098_ (.A(_09440_),
    .ZN(_09441_));
 OAI21_X1 _19099_ (.A(_08609_),
    .B1(_08697_),
    .B2(_08568_),
    .ZN(_09442_));
 NAND3_X1 _19100_ (.A1(_08655_),
    .A2(_08641_),
    .A3(_08642_),
    .ZN(_09443_));
 AND4_X1 _19101_ (.A1(_09439_),
    .A2(_09441_),
    .A3(_09442_),
    .A4(_09443_),
    .ZN(_09444_));
 AND4_X1 _19102_ (.A1(_09429_),
    .A2(_09435_),
    .A3(_09438_),
    .A4(_09444_),
    .ZN(_09445_));
 NAND4_X1 _19103_ (.A1(_09393_),
    .A2(_09410_),
    .A3(_09428_),
    .A4(_09445_),
    .ZN(_09446_));
 NOR2_X2 _19104_ (.A1(_09446_),
    .A2(_08696_),
    .ZN(_09447_));
 XNOR2_X2 _19105_ (.A(_09372_),
    .B(_09447_),
    .ZN(_09448_));
 XNOR2_X1 _19106_ (.A(_09448_),
    .B(_08814_),
    .ZN(_09449_));
 XNOR2_X1 _19107_ (.A(_09259_),
    .B(_09449_),
    .ZN(_09450_));
 INV_X1 _19108_ (.A(_17078_),
    .ZN(_09451_));
 BUF_X2 _19109_ (.A(_09451_),
    .Z(_09452_));
 XNOR2_X1 _19110_ (.A(_09450_),
    .B(_09452_),
    .ZN(_09453_));
 MUX2_X1 _19111_ (.A(_09042_),
    .B(_09453_),
    .S(_09040_),
    .Z(_00725_));
 XOR2_X1 _19112_ (.A(_17089_),
    .B(_16985_),
    .Z(_09454_));
 AOI211_X1 _19113_ (.A(_06842_),
    .B(_08492_),
    .C1(_08459_),
    .C2(_07161_),
    .ZN(_09455_));
 BUF_X2 _19114_ (.A(_09263_),
    .Z(_09456_));
 NAND2_X1 _19115_ (.A1(_08491_),
    .A2(_09456_),
    .ZN(_09457_));
 OAI211_X1 _19116_ (.A(_09275_),
    .B(_09457_),
    .C1(_09349_),
    .C2(_08492_),
    .ZN(_09458_));
 AND3_X1 _19117_ (.A1(_08167_),
    .A2(_08200_),
    .A3(_07543_),
    .ZN(_09459_));
 NOR3_X1 _19118_ (.A1(_09455_),
    .A2(_09458_),
    .A3(_09459_),
    .ZN(_09460_));
 NAND2_X1 _19119_ (.A1(_07466_),
    .A2(_08451_),
    .ZN(_09461_));
 OAI21_X1 _19120_ (.A(_09461_),
    .B1(_09346_),
    .B2(_07707_),
    .ZN(_09462_));
 NAND3_X1 _19121_ (.A1(_09330_),
    .A2(_08211_),
    .A3(_06699_),
    .ZN(_09463_));
 OAI21_X1 _19122_ (.A(_09463_),
    .B1(_09346_),
    .B2(_09287_),
    .ZN(_09464_));
 AND3_X1 _19123_ (.A1(_08211_),
    .A2(_07183_),
    .A3(_06699_),
    .ZN(_09465_));
 AND2_X1 _19124_ (.A1(_07455_),
    .A2(_07367_),
    .ZN(_09466_));
 NOR4_X1 _19125_ (.A1(_09462_),
    .A2(_09464_),
    .A3(_09465_),
    .A4(_09466_),
    .ZN(_09467_));
 INV_X2 _19126_ (.A(_06831_),
    .ZN(_09468_));
 AOI211_X1 _19127_ (.A(_07128_),
    .B(_09468_),
    .C1(_06754_),
    .C2(_08091_),
    .ZN(_09469_));
 AOI21_X1 _19128_ (.A(_09468_),
    .B1(_08327_),
    .B2(_09310_),
    .ZN(_09470_));
 AND4_X1 _19129_ (.A1(_06853_),
    .A2(_06809_),
    .A3(_07356_),
    .A4(_07554_),
    .ZN(_09471_));
 NOR4_X1 _19130_ (.A1(_09469_),
    .A2(_06897_),
    .A3(_09470_),
    .A4(_09471_),
    .ZN(_09472_));
 AND2_X1 _19131_ (.A1(_09352_),
    .A2(_07378_),
    .ZN(_09473_));
 AND2_X1 _19132_ (.A1(_09351_),
    .A2(_06765_),
    .ZN(_09474_));
 AND3_X1 _19133_ (.A1(_07937_),
    .A2(_07992_),
    .A3(_08211_),
    .ZN(_09475_));
 NOR4_X1 _19134_ (.A1(_09473_),
    .A2(_09357_),
    .A3(_09474_),
    .A4(_09475_),
    .ZN(_09476_));
 AND2_X1 _19135_ (.A1(_07631_),
    .A2(_09327_),
    .ZN(_09477_));
 OAI21_X1 _19136_ (.A(_09362_),
    .B1(_07641_),
    .B2(_07510_),
    .ZN(_09478_));
 AOI211_X1 _19137_ (.A(_09477_),
    .B(_09478_),
    .C1(_08467_),
    .C2(_07631_),
    .ZN(_09479_));
 AND4_X1 _19138_ (.A1(_09467_),
    .A2(_09472_),
    .A3(_09476_),
    .A4(_09479_),
    .ZN(_09480_));
 OAI21_X1 _19139_ (.A(_07576_),
    .B1(_09289_),
    .B2(_08455_),
    .ZN(_09481_));
 NAND3_X1 _19140_ (.A1(_08384_),
    .A2(_07576_),
    .A3(_09325_),
    .ZN(_09482_));
 OAI211_X1 _19141_ (.A(_09481_),
    .B(_09482_),
    .C1(_09310_),
    .C2(_09261_),
    .ZN(_09483_));
 INV_X1 _19142_ (.A(_07378_),
    .ZN(_09484_));
 AOI21_X1 _19143_ (.A(_07293_),
    .B1(_09277_),
    .B2(_09484_),
    .ZN(_09485_));
 AND2_X1 _19144_ (.A1(_08167_),
    .A2(_07007_),
    .ZN(_09486_));
 AND3_X1 _19145_ (.A1(_07861_),
    .A2(_08431_),
    .A3(_07007_),
    .ZN(_09487_));
 NOR4_X1 _19146_ (.A1(_09483_),
    .A2(_09485_),
    .A3(_09486_),
    .A4(_09487_),
    .ZN(_09488_));
 OAI211_X1 _19147_ (.A(_07238_),
    .B(_08069_),
    .C1(_06754_),
    .C2(_08091_),
    .ZN(_09489_));
 NAND2_X1 _19148_ (.A1(_09313_),
    .A2(_07238_),
    .ZN(_09490_));
 NAND2_X1 _19149_ (.A1(_09489_),
    .A2(_09490_),
    .ZN(_09491_));
 AOI21_X1 _19150_ (.A(_08481_),
    .B1(_07510_),
    .B2(_09310_),
    .ZN(_09492_));
 AOI211_X1 _19151_ (.A(_09491_),
    .B(_09492_),
    .C1(_07249_),
    .C2(_06776_),
    .ZN(_09493_));
 AND4_X1 _19152_ (.A1(_09460_),
    .A2(_09480_),
    .A3(_09488_),
    .A4(_09493_),
    .ZN(_09494_));
 OAI21_X1 _19153_ (.A(_07411_),
    .B1(_07806_),
    .B2(_08455_),
    .ZN(_09495_));
 NAND4_X1 _19154_ (.A1(_07554_),
    .A2(_08478_),
    .A3(_08463_),
    .A4(_06930_),
    .ZN(_09496_));
 NAND4_X1 _19155_ (.A1(_07400_),
    .A2(_07194_),
    .A3(_07850_),
    .A4(_08431_),
    .ZN(_09497_));
 AND3_X1 _19156_ (.A1(_09495_),
    .A2(_09496_),
    .A3(_09497_),
    .ZN(_09498_));
 AND2_X1 _19157_ (.A1(_08145_),
    .A2(_08451_),
    .ZN(_09499_));
 AND2_X1 _19158_ (.A1(_08145_),
    .A2(_08308_),
    .ZN(_09500_));
 AND3_X1 _19159_ (.A1(_08455_),
    .A2(_07992_),
    .A3(_07062_),
    .ZN(_09501_));
 OR4_X1 _19160_ (.A1(_09499_),
    .A2(_09328_),
    .A3(_09500_),
    .A4(_09501_),
    .ZN(_09502_));
 OAI21_X1 _19161_ (.A(_07084_),
    .B1(_07981_),
    .B2(_08467_),
    .ZN(_09503_));
 AND2_X1 _19162_ (.A1(_07084_),
    .A2(_07532_),
    .ZN(_09504_));
 INV_X1 _19163_ (.A(_09504_),
    .ZN(_09505_));
 NAND2_X1 _19164_ (.A1(_08308_),
    .A2(_07084_),
    .ZN(_09506_));
 NAND2_X1 _19165_ (.A1(_07084_),
    .A2(_09321_),
    .ZN(_09507_));
 NAND4_X1 _19166_ (.A1(_09503_),
    .A2(_09505_),
    .A3(_09506_),
    .A4(_09507_),
    .ZN(_09508_));
 OAI21_X1 _19167_ (.A(_07893_),
    .B1(_09327_),
    .B2(_09263_),
    .ZN(_09509_));
 OAI21_X1 _19168_ (.A(_09509_),
    .B1(_08494_),
    .B2(_09311_),
    .ZN(_09510_));
 AND2_X1 _19169_ (.A1(_09313_),
    .A2(_07674_),
    .ZN(_09511_));
 INV_X1 _19170_ (.A(_09511_),
    .ZN(_09512_));
 AND2_X1 _19171_ (.A1(_09330_),
    .A2(_07674_),
    .ZN(_09513_));
 INV_X1 _19172_ (.A(_09513_),
    .ZN(_09514_));
 AND2_X1 _19173_ (.A1(_07674_),
    .A2(_08451_),
    .ZN(_09515_));
 INV_X1 _19174_ (.A(_09515_),
    .ZN(_09516_));
 NAND4_X1 _19175_ (.A1(_09512_),
    .A2(_09514_),
    .A3(_09516_),
    .A4(_08499_),
    .ZN(_09517_));
 NOR4_X1 _19176_ (.A1(_09502_),
    .A2(_09508_),
    .A3(_09510_),
    .A4(_09517_),
    .ZN(_09518_));
 OAI21_X1 _19177_ (.A(_08025_),
    .B1(_09330_),
    .B2(_07948_),
    .ZN(_09519_));
 OAI21_X1 _19178_ (.A(_08025_),
    .B1(_07795_),
    .B2(_08451_),
    .ZN(_09520_));
 OAI211_X1 _19179_ (.A(_09519_),
    .B(_09520_),
    .C1(_09484_),
    .C2(_09292_),
    .ZN(_09521_));
 NAND2_X1 _19180_ (.A1(_09324_),
    .A2(_06721_),
    .ZN(_09522_));
 NAND4_X1 _19181_ (.A1(_07150_),
    .A2(_08069_),
    .A3(_06699_),
    .A4(_08463_),
    .ZN(_09523_));
 NAND2_X1 _19182_ (.A1(_09522_),
    .A2(_09523_),
    .ZN(_09524_));
 NAND2_X1 _19183_ (.A1(_08473_),
    .A2(_06732_),
    .ZN(_09525_));
 OAI22_X1 _19184_ (.A1(_09525_),
    .A2(_07598_),
    .B1(_07510_),
    .B2(_07488_),
    .ZN(_09526_));
 NOR3_X1 _19185_ (.A1(_09521_),
    .A2(_09524_),
    .A3(_09526_),
    .ZN(_09527_));
 OAI21_X1 _19186_ (.A(_07839_),
    .B1(_08167_),
    .B2(_06952_),
    .ZN(_09528_));
 OAI211_X1 _19187_ (.A(_07839_),
    .B(_08069_),
    .C1(_06930_),
    .C2(_07161_),
    .ZN(_09529_));
 NAND2_X1 _19188_ (.A1(_07839_),
    .A2(_08384_),
    .ZN(_09530_));
 NAND4_X1 _19189_ (.A1(_06974_),
    .A2(_07598_),
    .A3(_08233_),
    .A4(_08463_),
    .ZN(_09531_));
 AND4_X1 _19190_ (.A1(_09528_),
    .A2(_09529_),
    .A3(_09530_),
    .A4(_09531_),
    .ZN(_09532_));
 AND4_X1 _19191_ (.A1(_09498_),
    .A2(_09518_),
    .A3(_09527_),
    .A4(_09532_),
    .ZN(_09533_));
 NAND2_X2 _19192_ (.A1(_09494_),
    .A2(_09533_),
    .ZN(_09534_));
 AND2_X1 _19193_ (.A1(_08585_),
    .A2(_08684_),
    .ZN(_09535_));
 AND2_X1 _19194_ (.A1(_08584_),
    .A2(_08620_),
    .ZN(_09536_));
 AND2_X1 _19195_ (.A1(_08584_),
    .A2(_08665_),
    .ZN(_09537_));
 OR3_X1 _19196_ (.A1(_09535_),
    .A2(_09536_),
    .A3(_09537_),
    .ZN(_09538_));
 AND2_X1 _19197_ (.A1(_08585_),
    .A2(_08573_),
    .ZN(_09539_));
 AND3_X1 _19198_ (.A1(_08764_),
    .A2(_08540_),
    .A3(_08581_),
    .ZN(_09540_));
 AND2_X1 _19199_ (.A1(_08585_),
    .A2(_08578_),
    .ZN(_09541_));
 NOR4_X1 _19200_ (.A1(_09538_),
    .A2(_09539_),
    .A3(_09540_),
    .A4(_09541_),
    .ZN(_09542_));
 AND2_X1 _19201_ (.A1(_08588_),
    .A2(_08590_),
    .ZN(_09543_));
 OAI21_X1 _19202_ (.A(_08636_),
    .B1(_09543_),
    .B2(_08724_),
    .ZN(_09544_));
 OAI21_X1 _19203_ (.A(_08636_),
    .B1(_08715_),
    .B2(_08682_),
    .ZN(_09545_));
 AND3_X1 _19204_ (.A1(_09542_),
    .A2(_09544_),
    .A3(_09545_),
    .ZN(_09546_));
 INV_X1 _19205_ (.A(_08536_),
    .ZN(_09547_));
 AND2_X1 _19206_ (.A1(_08774_),
    .A2(_08590_),
    .ZN(_09548_));
 INV_X1 _19207_ (.A(_09548_),
    .ZN(_09549_));
 AOI21_X1 _19208_ (.A(_08767_),
    .B1(_09547_),
    .B2(_09549_),
    .ZN(_09550_));
 AOI21_X1 _19209_ (.A(_08558_),
    .B1(_08710_),
    .B2(_08802_),
    .ZN(_09551_));
 NAND2_X1 _19210_ (.A1(_08565_),
    .A2(_08689_),
    .ZN(_09552_));
 NAND2_X1 _19211_ (.A1(_08565_),
    .A2(_08704_),
    .ZN(_09553_));
 OAI211_X1 _19212_ (.A(_09552_),
    .B(_09553_),
    .C1(_08767_),
    .C2(_09417_),
    .ZN(_09554_));
 NOR4_X1 _19213_ (.A1(_09550_),
    .A2(_08555_),
    .A3(_09551_),
    .A4(_09554_),
    .ZN(_09555_));
 OAI21_X1 _19214_ (.A(_08629_),
    .B1(_08704_),
    .B2(_08594_),
    .ZN(_09556_));
 OAI21_X1 _19215_ (.A(_08629_),
    .B1(_08764_),
    .B2(_08607_),
    .ZN(_09557_));
 OAI21_X1 _19216_ (.A(_08664_),
    .B1(_08704_),
    .B2(_08553_),
    .ZN(_09558_));
 OAI21_X1 _19217_ (.A(_08664_),
    .B1(_08764_),
    .B2(_08682_),
    .ZN(_09559_));
 AND4_X1 _19218_ (.A1(_09556_),
    .A2(_09557_),
    .A3(_09558_),
    .A4(_09559_),
    .ZN(_09560_));
 NAND3_X1 _19219_ (.A1(_08797_),
    .A2(_08657_),
    .A3(_08539_),
    .ZN(_09561_));
 AND2_X1 _19220_ (.A1(_08620_),
    .A2(_08599_),
    .ZN(_09562_));
 AND3_X1 _19221_ (.A1(_08672_),
    .A2(_08598_),
    .A3(_08587_),
    .ZN(_09563_));
 MUX2_X1 _19222_ (.A(_08567_),
    .B(_08631_),
    .S(_08534_),
    .Z(_09564_));
 AOI211_X1 _19223_ (.A(_09562_),
    .B(_09563_),
    .C1(_08622_),
    .C2(_09564_),
    .ZN(_09565_));
 OAI21_X1 _19224_ (.A(_08542_),
    .B1(_08714_),
    .B2(_08553_),
    .ZN(_09566_));
 OAI211_X1 _19225_ (.A(_08542_),
    .B(_08733_),
    .C1(_09382_),
    .C2(_08574_),
    .ZN(_09567_));
 AND4_X1 _19226_ (.A1(_09561_),
    .A2(_09565_),
    .A3(_09566_),
    .A4(_09567_),
    .ZN(_09568_));
 NAND4_X1 _19227_ (.A1(_09546_),
    .A2(_09555_),
    .A3(_09560_),
    .A4(_09568_),
    .ZN(_09569_));
 OAI21_X1 _19228_ (.A(_08650_),
    .B1(_08621_),
    .B2(_08685_),
    .ZN(_09570_));
 AND2_X1 _19229_ (.A1(_08604_),
    .A2(_08600_),
    .ZN(_09571_));
 INV_X1 _19230_ (.A(_08604_),
    .ZN(_09572_));
 AOI21_X1 _19231_ (.A(_09572_),
    .B1(_08693_),
    .B2(_08802_),
    .ZN(_09573_));
 AOI211_X1 _19232_ (.A(_09571_),
    .B(_09573_),
    .C1(_08605_),
    .C2(_08797_),
    .ZN(_09574_));
 OAI21_X1 _19233_ (.A(_08649_),
    .B1(_08553_),
    .B2(_08724_),
    .ZN(_09575_));
 OAI211_X1 _19234_ (.A(_08650_),
    .B(_16706_),
    .C1(_08574_),
    .C2(_08515_),
    .ZN(_09576_));
 AND4_X1 _19235_ (.A1(_09570_),
    .A2(_09574_),
    .A3(_09575_),
    .A4(_09576_),
    .ZN(_09577_));
 INV_X1 _19236_ (.A(_08611_),
    .ZN(_09578_));
 OAI211_X1 _19237_ (.A(_09441_),
    .B(_08757_),
    .C1(_08754_),
    .C2(_09578_),
    .ZN(_09579_));
 AOI21_X1 _19238_ (.A(_08752_),
    .B1(_09549_),
    .B2(_09390_),
    .ZN(_09580_));
 INV_X1 _19239_ (.A(_08620_),
    .ZN(_09581_));
 AOI21_X1 _19240_ (.A(_08752_),
    .B1(_08711_),
    .B2(_09581_),
    .ZN(_09582_));
 NAND3_X1 _19241_ (.A1(_08578_),
    .A2(_08641_),
    .A3(_08642_),
    .ZN(_09583_));
 NAND4_X1 _19242_ (.A1(_08641_),
    .A2(_08631_),
    .A3(_08618_),
    .A4(_08521_),
    .ZN(_09584_));
 INV_X1 _19243_ (.A(_08661_),
    .ZN(_09585_));
 OAI211_X1 _19244_ (.A(_09583_),
    .B(_09584_),
    .C1(_08754_),
    .C2(_09585_),
    .ZN(_09586_));
 NOR4_X1 _19245_ (.A1(_09579_),
    .A2(_09580_),
    .A3(_09582_),
    .A4(_09586_),
    .ZN(_09587_));
 OAI21_X1 _19246_ (.A(_08677_),
    .B1(_08746_),
    .B2(_08732_),
    .ZN(_09588_));
 OAI21_X1 _19247_ (.A(_08523_),
    .B1(_08708_),
    .B2(_08682_),
    .ZN(_09589_));
 OAI21_X1 _19248_ (.A(_08523_),
    .B1(_08681_),
    .B2(_08685_),
    .ZN(_09590_));
 AND4_X1 _19249_ (.A1(_08726_),
    .A2(_09588_),
    .A3(_09589_),
    .A4(_09590_),
    .ZN(_09591_));
 OAI21_X1 _19250_ (.A(_08703_),
    .B1(_08689_),
    .B2(_08601_),
    .ZN(_09592_));
 NAND3_X1 _19251_ (.A1(_08667_),
    .A2(_08703_),
    .A3(_08590_),
    .ZN(_09593_));
 OAI21_X1 _19252_ (.A(_08703_),
    .B1(_08640_),
    .B2(_08607_),
    .ZN(_09594_));
 NAND4_X1 _19253_ (.A1(_09592_),
    .A2(_09593_),
    .A3(_09594_),
    .A4(_09376_),
    .ZN(_09595_));
 OAI211_X1 _19254_ (.A(_08592_),
    .B(_08733_),
    .C1(_09382_),
    .C2(_08794_),
    .ZN(_09596_));
 NAND2_X1 _19255_ (.A1(_08698_),
    .A2(_08592_),
    .ZN(_09597_));
 NAND2_X1 _19256_ (.A1(_09596_),
    .A2(_09597_),
    .ZN(_09598_));
 INV_X1 _19257_ (.A(_08601_),
    .ZN(_09599_));
 AOI21_X1 _19258_ (.A(_08529_),
    .B1(_08669_),
    .B2(_09599_),
    .ZN(_09600_));
 NOR3_X1 _19259_ (.A1(_09595_),
    .A2(_09598_),
    .A3(_09600_),
    .ZN(_09601_));
 NAND4_X1 _19260_ (.A1(_09577_),
    .A2(_09587_),
    .A3(_09591_),
    .A4(_09601_),
    .ZN(_09602_));
 NOR2_X2 _19261_ (.A1(_09569_),
    .A2(_09602_),
    .ZN(_09603_));
 XNOR2_X1 _19262_ (.A(_09534_),
    .B(_09603_),
    .ZN(_09604_));
 NAND2_X1 _19263_ (.A1(_05064_),
    .A2(_05896_),
    .ZN(_09605_));
 NAND2_X1 _19264_ (.A1(_05599_),
    .A2(_06017_),
    .ZN(_09606_));
 NAND3_X1 _19265_ (.A1(_06017_),
    .A2(_04329_),
    .A3(_04658_),
    .ZN(_09607_));
 INV_X1 _19266_ (.A(_05962_),
    .ZN(_09608_));
 OAI211_X1 _19267_ (.A(_09606_),
    .B(_09607_),
    .C1(_09248_),
    .C2(_09608_),
    .ZN(_09609_));
 AOI211_X1 _19268_ (.A(_09244_),
    .B(_09609_),
    .C1(_09246_),
    .C2(_05929_),
    .ZN(_09610_));
 NAND3_X1 _19269_ (.A1(_06468_),
    .A2(_05907_),
    .A3(_04899_),
    .ZN(_09611_));
 NOR2_X2 _19270_ (.A1(_04910_),
    .A2(_04253_),
    .ZN(_09612_));
 NAND2_X1 _19271_ (.A1(_09612_),
    .A2(_05907_),
    .ZN(_09613_));
 AND4_X1 _19272_ (.A1(_09605_),
    .A2(_09610_),
    .A3(_09611_),
    .A4(_09613_),
    .ZN(_09614_));
 AND2_X1 _19273_ (.A1(_05313_),
    .A2(_04658_),
    .ZN(_09615_));
 NAND3_X1 _19274_ (.A1(_09615_),
    .A2(_09158_),
    .A3(_05874_),
    .ZN(_09616_));
 NAND2_X1 _19275_ (.A1(_05632_),
    .A2(_06490_),
    .ZN(_09617_));
 NAND2_X1 _19276_ (.A1(_05632_),
    .A2(_05159_),
    .ZN(_09618_));
 NAND4_X1 _19277_ (.A1(_05621_),
    .A2(_09616_),
    .A3(_09617_),
    .A4(_09618_),
    .ZN(_09619_));
 NAND3_X1 _19278_ (.A1(_05064_),
    .A2(_05687_),
    .A3(_05874_),
    .ZN(_09620_));
 NAND2_X1 _19279_ (.A1(_05632_),
    .A2(_04778_),
    .ZN(_09621_));
 OAI221_X1 _19280_ (.A(_09620_),
    .B1(_05654_),
    .B2(_05434_),
    .C1(_05192_),
    .C2(_09621_),
    .ZN(_09622_));
 BUF_X2 _19281_ (.A(_09149_),
    .Z(_09623_));
 OAI21_X1 _19282_ (.A(_05775_),
    .B1(_09623_),
    .B2(_05082_),
    .ZN(_09624_));
 NAND2_X1 _19283_ (.A1(_05599_),
    .A2(_05775_),
    .ZN(_09625_));
 NAND2_X1 _19284_ (.A1(_09624_),
    .A2(_09625_),
    .ZN(_09626_));
 OAI211_X1 _19285_ (.A(_05775_),
    .B(_04713_),
    .C1(_05313_),
    .C2(_04735_),
    .ZN(_09627_));
 NAND3_X1 _19286_ (.A1(_05775_),
    .A2(_05137_),
    .A3(_04713_),
    .ZN(_09628_));
 OAI211_X1 _19287_ (.A(_09627_),
    .B(_09628_),
    .C1(_05434_),
    .C2(_09238_),
    .ZN(_09629_));
 NOR4_X1 _19288_ (.A1(_09619_),
    .A2(_09622_),
    .A3(_09626_),
    .A4(_09629_),
    .ZN(_09630_));
 NOR2_X1 _19289_ (.A1(_06402_),
    .A2(_04253_),
    .ZN(_09631_));
 NAND2_X1 _19290_ (.A1(_05511_),
    .A2(_09631_),
    .ZN(_09632_));
 AND2_X1 _19291_ (.A1(_05214_),
    .A2(_04625_),
    .ZN(_09633_));
 AND3_X1 _19292_ (.A1(_04548_),
    .A2(_05687_),
    .A3(_05110_),
    .ZN(_09634_));
 NOR4_X1 _19293_ (.A1(_05236_),
    .A2(_09633_),
    .A3(_09161_),
    .A4(_09634_),
    .ZN(_09635_));
 OAI21_X1 _19294_ (.A(_05511_),
    .B1(_05064_),
    .B2(_04307_),
    .ZN(_09636_));
 OAI211_X1 _19295_ (.A(_05511_),
    .B(_16754_),
    .C1(_04959_),
    .C2(_04220_),
    .ZN(_09637_));
 AND4_X1 _19296_ (.A1(_09632_),
    .A2(_09635_),
    .A3(_09636_),
    .A4(_09637_),
    .ZN(_09638_));
 AND2_X1 _19297_ (.A1(_04921_),
    .A2(_04899_),
    .ZN(_09639_));
 OAI21_X1 _19298_ (.A(_05291_),
    .B1(_09639_),
    .B2(_05599_),
    .ZN(_09640_));
 NAND2_X1 _19299_ (.A1(_04263_),
    .A2(_05258_),
    .ZN(_09641_));
 AND2_X1 _19300_ (.A1(_05258_),
    .A2(_04340_),
    .ZN(_09642_));
 INV_X1 _19301_ (.A(_09642_),
    .ZN(_09643_));
 NAND4_X1 _19302_ (.A1(_09640_),
    .A2(_09179_),
    .A3(_09641_),
    .A4(_09643_),
    .ZN(_09644_));
 AOI211_X1 _19303_ (.A(_05357_),
    .B(_05423_),
    .C1(_05137_),
    .C2(_04680_),
    .ZN(_09645_));
 OAI21_X1 _19304_ (.A(_05401_),
    .B1(_04395_),
    .B2(_05478_),
    .ZN(_09646_));
 NAND4_X1 _19305_ (.A1(_05368_),
    .A2(_04669_),
    .A3(_05324_),
    .A4(_04833_),
    .ZN(_09647_));
 OAI211_X1 _19306_ (.A(_09646_),
    .B(_09647_),
    .C1(_05423_),
    .C2(_04526_),
    .ZN(_09648_));
 NOR4_X1 _19307_ (.A1(_09644_),
    .A2(_09645_),
    .A3(_05467_),
    .A4(_09648_),
    .ZN(_09649_));
 NAND4_X1 _19308_ (.A1(_09614_),
    .A2(_09630_),
    .A3(_09638_),
    .A4(_09649_),
    .ZN(_09650_));
 NAND2_X1 _19309_ (.A1(_06160_),
    .A2(_04636_),
    .ZN(_09651_));
 AND3_X1 _19310_ (.A1(_06413_),
    .A2(_06236_),
    .A3(_06270_),
    .ZN(_09652_));
 AND2_X1 _19311_ (.A1(_09612_),
    .A2(_06270_),
    .ZN(_09653_));
 AND2_X1 _19312_ (.A1(_05064_),
    .A2(_06270_),
    .ZN(_09654_));
 NOR4_X1 _19313_ (.A1(_09652_),
    .A2(_09653_),
    .A3(_09654_),
    .A4(_09216_),
    .ZN(_09655_));
 OAI21_X1 _19314_ (.A(_06160_),
    .B1(_04263_),
    .B2(_05017_),
    .ZN(_09656_));
 OAI21_X1 _19315_ (.A(_06160_),
    .B1(_04537_),
    .B2(_04559_),
    .ZN(_09657_));
 AND4_X1 _19316_ (.A1(_09651_),
    .A2(_09655_),
    .A3(_09656_),
    .A4(_09657_),
    .ZN(_09658_));
 NAND2_X1 _19317_ (.A1(_04888_),
    .A2(_05017_),
    .ZN(_09659_));
 NAND2_X1 _19318_ (.A1(_04888_),
    .A2(_09623_),
    .ZN(_09660_));
 NAND2_X1 _19319_ (.A1(_04888_),
    .A2(_04537_),
    .ZN(_09661_));
 NAND4_X1 _19320_ (.A1(_04877_),
    .A2(_09659_),
    .A3(_09660_),
    .A4(_09661_),
    .ZN(_09662_));
 AND2_X1 _19321_ (.A1(_04209_),
    .A2(_09149_),
    .ZN(_09663_));
 OR2_X1 _19322_ (.A1(_04406_),
    .A2(_09663_),
    .ZN(_09664_));
 AND2_X1 _19323_ (.A1(_06138_),
    .A2(_04209_),
    .ZN(_09665_));
 NAND2_X1 _19324_ (.A1(_04209_),
    .A2(_05120_),
    .ZN(_09666_));
 OAI211_X1 _19325_ (.A(_09666_),
    .B(_04351_),
    .C1(_04318_),
    .C2(_05192_),
    .ZN(_09667_));
 NOR4_X1 _19326_ (.A1(_09662_),
    .A2(_09664_),
    .A3(_09665_),
    .A4(_09667_),
    .ZN(_09668_));
 OAI21_X1 _19327_ (.A(_04614_),
    .B1(_09178_),
    .B2(_05676_),
    .ZN(_09669_));
 OAI21_X1 _19328_ (.A(_05045_),
    .B1(_09178_),
    .B2(_05017_),
    .ZN(_09670_));
 OAI21_X1 _19329_ (.A(_05045_),
    .B1(_05599_),
    .B2(_05962_),
    .ZN(_09671_));
 OAI21_X1 _19330_ (.A(_04614_),
    .B1(_05599_),
    .B2(_05159_),
    .ZN(_09672_));
 AND4_X1 _19331_ (.A1(_09669_),
    .A2(_09670_),
    .A3(_09671_),
    .A4(_09672_),
    .ZN(_09673_));
 OAI21_X1 _19332_ (.A(_06556_),
    .B1(_06238_),
    .B2(_04778_),
    .ZN(_09674_));
 OAI211_X1 _19333_ (.A(_06391_),
    .B(_04658_),
    .C1(_04242_),
    .C2(_05116_),
    .ZN(_09675_));
 NAND4_X1 _19334_ (.A1(_04472_),
    .A2(_04329_),
    .A3(_04384_),
    .A4(_06149_),
    .ZN(_09676_));
 AND2_X1 _19335_ (.A1(_09675_),
    .A2(_09676_),
    .ZN(_09677_));
 OAI21_X1 _19336_ (.A(_06556_),
    .B1(_06116_),
    .B2(_05962_),
    .ZN(_09678_));
 NAND2_X1 _19337_ (.A1(_06391_),
    .A2(_04296_),
    .ZN(_09679_));
 NAND2_X1 _19338_ (.A1(_06391_),
    .A2(_05064_),
    .ZN(_09680_));
 NAND2_X1 _19339_ (.A1(_06391_),
    .A2(_09631_),
    .ZN(_09681_));
 AND3_X1 _19340_ (.A1(_09679_),
    .A2(_09680_),
    .A3(_09681_),
    .ZN(_09682_));
 AND4_X1 _19341_ (.A1(_09674_),
    .A2(_09677_),
    .A3(_09678_),
    .A4(_09682_),
    .ZN(_09683_));
 NAND4_X1 _19342_ (.A1(_09658_),
    .A2(_09668_),
    .A3(_09673_),
    .A4(_09683_),
    .ZN(_09684_));
 NOR2_X2 _19343_ (.A1(_09650_),
    .A2(_09684_),
    .ZN(_09685_));
 XNOR2_X1 _19344_ (.A(_09604_),
    .B(_09685_),
    .ZN(_09686_));
 AND2_X1 _19345_ (.A1(_09062_),
    .A2(_08865_),
    .ZN(_09687_));
 AND3_X1 _19346_ (.A1(_08828_),
    .A2(_09107_),
    .A3(_08867_),
    .ZN(_09688_));
 NOR2_X1 _19347_ (.A1(_09687_),
    .A2(_09688_),
    .ZN(_09689_));
 AND2_X1 _19348_ (.A1(_08877_),
    .A2(_08822_),
    .ZN(_09690_));
 OAI21_X1 _19349_ (.A(_09106_),
    .B1(_08853_),
    .B2(_09690_),
    .ZN(_09691_));
 NAND3_X1 _19350_ (.A1(_09008_),
    .A2(_08844_),
    .A3(_08915_),
    .ZN(_09692_));
 NAND2_X1 _19351_ (.A1(_08906_),
    .A2(_09122_),
    .ZN(_09693_));
 NAND4_X1 _19352_ (.A1(_09689_),
    .A2(_09691_),
    .A3(_09692_),
    .A4(_09693_),
    .ZN(_09694_));
 NAND2_X1 _19353_ (.A1(_08986_),
    .A2(_08952_),
    .ZN(_09695_));
 NAND2_X1 _19354_ (.A1(_08987_),
    .A2(_08952_),
    .ZN(_09696_));
 NAND3_X1 _19355_ (.A1(_08889_),
    .A2(_08833_),
    .A3(_08950_),
    .ZN(_09697_));
 NAND3_X1 _19356_ (.A1(_09695_),
    .A2(_09696_),
    .A3(_09697_),
    .ZN(_09698_));
 AND2_X1 _19357_ (.A1(_09025_),
    .A2(_08915_),
    .ZN(_09699_));
 AND2_X1 _19358_ (.A1(_08976_),
    .A2(_08850_),
    .ZN(_09700_));
 OR3_X1 _19359_ (.A1(_09698_),
    .A2(_09699_),
    .A3(_09700_),
    .ZN(_09701_));
 NOR4_X1 _19360_ (.A1(_09694_),
    .A2(_09701_),
    .A3(_08920_),
    .A4(_09112_),
    .ZN(_09702_));
 NAND2_X1 _19361_ (.A1(_09021_),
    .A2(_08847_),
    .ZN(_09703_));
 AND3_X1 _19362_ (.A1(_08954_),
    .A2(_08913_),
    .A3(_08950_),
    .ZN(_09704_));
 AND2_X1 _19363_ (.A1(_09025_),
    .A2(_08942_),
    .ZN(_09705_));
 AND3_X1 _19364_ (.A1(_09093_),
    .A2(_08878_),
    .A3(_08957_),
    .ZN(_09706_));
 NOR4_X1 _19365_ (.A1(_09043_),
    .A2(_09704_),
    .A3(_09705_),
    .A4(_09706_),
    .ZN(_09707_));
 NAND2_X1 _19366_ (.A1(_09062_),
    .A2(_08940_),
    .ZN(_09708_));
 AND3_X1 _19367_ (.A1(_08853_),
    .A2(_08952_),
    .A3(_08844_),
    .ZN(_09709_));
 BUF_X2 _19368_ (.A(_09014_),
    .Z(_09710_));
 AOI21_X1 _19369_ (.A(_09709_),
    .B1(_09075_),
    .B2(_09710_),
    .ZN(_09711_));
 AND4_X1 _19370_ (.A1(_09703_),
    .A2(_09707_),
    .A3(_09708_),
    .A4(_09711_),
    .ZN(_09712_));
 AND4_X1 _19371_ (.A1(_08868_),
    .A2(_09115_),
    .A3(_09003_),
    .A4(_08827_),
    .ZN(_09713_));
 NOR2_X1 _19372_ (.A1(_09103_),
    .A2(_09713_),
    .ZN(_09714_));
 OAI21_X1 _19373_ (.A(_09016_),
    .B1(_08818_),
    .B2(_08867_),
    .ZN(_09715_));
 OAI21_X1 _19374_ (.A(_08936_),
    .B1(_09011_),
    .B2(_09715_),
    .ZN(_09716_));
 OAI21_X1 _19375_ (.A(_09031_),
    .B1(_09095_),
    .B2(_09093_),
    .ZN(_09717_));
 OAI21_X1 _19376_ (.A(_09005_),
    .B1(_08938_),
    .B2(_08860_),
    .ZN(_09718_));
 AND4_X1 _19377_ (.A1(_09714_),
    .A2(_09716_),
    .A3(_09717_),
    .A4(_09718_),
    .ZN(_09719_));
 BUF_X2 _19378_ (.A(_08901_),
    .Z(_09720_));
 OAI21_X1 _19379_ (.A(_09720_),
    .B1(_08938_),
    .B2(_09050_),
    .ZN(_09721_));
 NAND2_X1 _19380_ (.A1(_08929_),
    .A2(_08903_),
    .ZN(_09722_));
 NAND3_X1 _19381_ (.A1(_08930_),
    .A2(_09003_),
    .A3(_08913_),
    .ZN(_09723_));
 NAND2_X1 _19382_ (.A1(_08954_),
    .A2(_09031_),
    .ZN(_09724_));
 AND3_X1 _19383_ (.A1(_09722_),
    .A2(_09723_),
    .A3(_09724_),
    .ZN(_09725_));
 OAI21_X1 _19384_ (.A(_08941_),
    .B1(_09095_),
    .B2(_08889_),
    .ZN(_09726_));
 OAI21_X1 _19385_ (.A(_09053_),
    .B1(_09017_),
    .B2(_09077_),
    .ZN(_09727_));
 AND4_X1 _19386_ (.A1(_09721_),
    .A2(_09725_),
    .A3(_09726_),
    .A4(_09727_),
    .ZN(_09728_));
 NAND4_X1 _19387_ (.A1(_09702_),
    .A2(_09712_),
    .A3(_09719_),
    .A4(_09728_),
    .ZN(_09729_));
 AND2_X1 _19388_ (.A1(_08828_),
    .A2(_08842_),
    .ZN(_09730_));
 INV_X1 _19389_ (.A(_09730_),
    .ZN(_09731_));
 AND4_X1 _19390_ (.A1(_08854_),
    .A2(_08962_),
    .A3(_08922_),
    .A4(_09731_),
    .ZN(_09732_));
 AND2_X1 _19391_ (.A1(_08940_),
    .A2(_08874_),
    .ZN(_09733_));
 AND2_X1 _19392_ (.A1(_08923_),
    .A2(_08994_),
    .ZN(_09734_));
 NOR4_X1 _19393_ (.A1(_08837_),
    .A2(_09733_),
    .A3(_09734_),
    .A4(_08891_),
    .ZN(_09735_));
 AOI22_X1 _19394_ (.A1(_08847_),
    .A2(_09690_),
    .B1(_09007_),
    .B2(_08904_),
    .ZN(_09736_));
 NAND2_X1 _19395_ (.A1(_08929_),
    .A2(_08904_),
    .ZN(_09737_));
 NAND3_X1 _19396_ (.A1(_09048_),
    .A2(_08886_),
    .A3(_09003_),
    .ZN(_09738_));
 AND3_X1 _19397_ (.A1(_09736_),
    .A2(_09737_),
    .A3(_09738_),
    .ZN(_09739_));
 AND2_X1 _19398_ (.A1(_09026_),
    .A2(_09118_),
    .ZN(_09740_));
 AND2_X1 _19399_ (.A1(_08828_),
    .A2(_08915_),
    .ZN(_09741_));
 NOR4_X1 _19400_ (.A1(_09740_),
    .A2(_09060_),
    .A3(_09072_),
    .A4(_09741_),
    .ZN(_09742_));
 AND4_X1 _19401_ (.A1(_09732_),
    .A2(_09735_),
    .A3(_09739_),
    .A4(_09742_),
    .ZN(_09743_));
 OAI21_X1 _19402_ (.A(_08888_),
    .B1(_09021_),
    .B2(_09093_),
    .ZN(_09744_));
 AND3_X1 _19403_ (.A1(_09744_),
    .A2(_09137_),
    .A3(_09135_),
    .ZN(_09745_));
 AND4_X1 _19404_ (.A1(_08973_),
    .A2(_09087_),
    .A3(_16794_),
    .A4(_09088_),
    .ZN(_09746_));
 AND2_X1 _19405_ (.A1(_08954_),
    .A2(_09087_),
    .ZN(_09747_));
 AND2_X1 _19406_ (.A1(_09053_),
    .A2(_09009_),
    .ZN(_09748_));
 NOR3_X1 _19407_ (.A1(_09746_),
    .A2(_09747_),
    .A3(_09748_),
    .ZN(_09749_));
 INV_X1 _19408_ (.A(_08972_),
    .ZN(_09750_));
 OR2_X1 _19409_ (.A1(_09010_),
    .A2(_09750_),
    .ZN(_09751_));
 AND2_X1 _19410_ (.A1(_09128_),
    .A2(_09129_),
    .ZN(_09752_));
 NOR3_X1 _19411_ (.A1(_08978_),
    .A2(_09752_),
    .A3(_08980_),
    .ZN(_09753_));
 AOI22_X1 _19412_ (.A1(_09075_),
    .A2(_09048_),
    .B1(_09008_),
    .B2(_08998_),
    .ZN(_09754_));
 AOI22_X1 _19413_ (.A1(_08843_),
    .A2(_09008_),
    .B1(_08994_),
    .B2(_08909_),
    .ZN(_09755_));
 AND4_X1 _19414_ (.A1(_09751_),
    .A2(_09753_),
    .A3(_09754_),
    .A4(_09755_),
    .ZN(_09756_));
 NAND4_X1 _19415_ (.A1(_09743_),
    .A2(_09745_),
    .A3(_09749_),
    .A4(_09756_),
    .ZN(_09757_));
 NOR2_X2 _19416_ (.A1(_09729_),
    .A2(_09757_),
    .ZN(_09758_));
 INV_X1 _19417_ (.A(_09758_),
    .ZN(_09759_));
 XNOR2_X1 _19418_ (.A(_09447_),
    .B(_09759_),
    .ZN(_09760_));
 XNOR2_X1 _19419_ (.A(_09686_),
    .B(_09760_),
    .ZN(_09761_));
 XNOR2_X1 _19420_ (.A(_09761_),
    .B(_17089_),
    .ZN(_09762_));
 MUX2_X1 _19421_ (.A(_09454_),
    .B(_09762_),
    .S(_09040_),
    .Z(_00726_));
 XOR2_X1 _19422_ (.A(_17092_),
    .B(_16996_),
    .Z(_09763_));
 OAI21_X1 _19423_ (.A(_08649_),
    .B1(_09548_),
    .B2(_08707_),
    .ZN(_09764_));
 NAND4_X1 _19424_ (.A1(_08580_),
    .A2(_08633_),
    .A3(_08614_),
    .A4(_08653_),
    .ZN(_09765_));
 AND3_X1 _19425_ (.A1(_09764_),
    .A2(_09575_),
    .A3(_09765_),
    .ZN(_09766_));
 AND3_X1 _19426_ (.A1(_08544_),
    .A2(_08539_),
    .A3(_08580_),
    .ZN(_09767_));
 OR2_X1 _19427_ (.A1(_09571_),
    .A2(_09767_),
    .ZN(_09768_));
 AND2_X1 _19428_ (.A1(_08746_),
    .A2(_08604_),
    .ZN(_09769_));
 AOI211_X1 _19429_ (.A(_09768_),
    .B(_09769_),
    .C1(_08637_),
    .C2(_08605_),
    .ZN(_09770_));
 AOI21_X1 _19430_ (.A(_08754_),
    .B1(_08710_),
    .B2(_08768_),
    .ZN(_09771_));
 NAND4_X1 _19431_ (.A1(_08580_),
    .A2(_08579_),
    .A3(_08521_),
    .A4(_08593_),
    .ZN(_09772_));
 NAND4_X1 _19432_ (.A1(_08580_),
    .A2(_08653_),
    .A3(_08614_),
    .A4(_08521_),
    .ZN(_09773_));
 OAI211_X1 _19433_ (.A(_09772_),
    .B(_09773_),
    .C1(_08754_),
    .C2(_09581_),
    .ZN(_09774_));
 AND3_X1 _19434_ (.A1(_08608_),
    .A2(_08535_),
    .A3(_08531_),
    .ZN(_09775_));
 NOR3_X1 _19435_ (.A1(_09771_),
    .A2(_09774_),
    .A3(_09775_),
    .ZN(_09776_));
 NAND2_X1 _19436_ (.A1(_08571_),
    .A2(_08519_),
    .ZN(_09777_));
 NAND2_X1 _19437_ (.A1(_08571_),
    .A2(_08758_),
    .ZN(_09778_));
 NAND2_X1 _19438_ (.A1(_09777_),
    .A2(_09778_),
    .ZN(_09779_));
 AND2_X1 _19439_ (.A1(_08572_),
    .A2(_08573_),
    .ZN(_09780_));
 AND2_X1 _19440_ (.A1(_08572_),
    .A2(_08764_),
    .ZN(_09781_));
 NOR4_X1 _19441_ (.A1(_09779_),
    .A2(_09780_),
    .A3(_09781_),
    .A4(_09436_),
    .ZN(_09782_));
 AND4_X1 _19442_ (.A1(_09766_),
    .A2(_09770_),
    .A3(_09776_),
    .A4(_09782_),
    .ZN(_09783_));
 NAND3_X1 _19443_ (.A1(_08646_),
    .A2(_08618_),
    .A3(_08637_),
    .ZN(_09784_));
 OAI211_X1 _19444_ (.A(_08646_),
    .B(_08733_),
    .C1(_09382_),
    .C2(_08794_),
    .ZN(_09785_));
 OAI211_X1 _19445_ (.A(_08646_),
    .B(_08615_),
    .C1(_08509_),
    .C2(_08653_),
    .ZN(_09786_));
 OAI21_X1 _19446_ (.A(_08646_),
    .B1(_08679_),
    .B2(_08601_),
    .ZN(_09787_));
 AND4_X1 _19447_ (.A1(_09784_),
    .A2(_09785_),
    .A3(_09786_),
    .A4(_09787_),
    .ZN(_09788_));
 OAI21_X1 _19448_ (.A(_08677_),
    .B1(_08594_),
    .B2(_08689_),
    .ZN(_09789_));
 OAI21_X1 _19449_ (.A(_08677_),
    .B1(_08714_),
    .B2(_08685_),
    .ZN(_09790_));
 OAI21_X1 _19450_ (.A(_08677_),
    .B1(_08510_),
    .B2(_08578_),
    .ZN(_09791_));
 OAI211_X1 _19451_ (.A(_08675_),
    .B(_08581_),
    .C1(_08640_),
    .C2(_08607_),
    .ZN(_09792_));
 AND4_X1 _19452_ (.A1(_09789_),
    .A2(_09790_),
    .A3(_09791_),
    .A4(_09792_),
    .ZN(_09793_));
 OAI21_X1 _19453_ (.A(_08703_),
    .B1(_08510_),
    .B2(_08606_),
    .ZN(_09794_));
 NAND4_X1 _19454_ (.A1(_08702_),
    .A2(_08535_),
    .A3(_08731_),
    .A4(_08615_),
    .ZN(_09795_));
 INV_X1 _19455_ (.A(_08689_),
    .ZN(_09796_));
 OAI211_X1 _19456_ (.A(_09794_),
    .B(_09795_),
    .C1(_09796_),
    .C2(_09373_),
    .ZN(_09797_));
 NAND4_X1 _19457_ (.A1(_08509_),
    .A2(_08675_),
    .A3(_08633_),
    .A4(_08593_),
    .ZN(_09798_));
 NAND4_X1 _19458_ (.A1(_08614_),
    .A2(_08633_),
    .A3(_08675_),
    .A4(_08653_),
    .ZN(_09799_));
 OAI211_X1 _19459_ (.A(_09798_),
    .B(_09799_),
    .C1(_08529_),
    .C2(_08557_),
    .ZN(_09800_));
 NAND2_X1 _19460_ (.A1(_08592_),
    .A2(_08797_),
    .ZN(_09801_));
 OAI21_X1 _19461_ (.A(_09801_),
    .B1(_08768_),
    .B2(_08529_),
    .ZN(_09802_));
 OAI21_X1 _19462_ (.A(_08514_),
    .B1(_08802_),
    .B2(_08529_),
    .ZN(_09803_));
 NOR4_X1 _19463_ (.A1(_09797_),
    .A2(_09800_),
    .A3(_09802_),
    .A4(_09803_),
    .ZN(_09804_));
 NAND4_X1 _19464_ (.A1(_09783_),
    .A2(_09788_),
    .A3(_09793_),
    .A4(_09804_),
    .ZN(_09805_));
 INV_X1 _19465_ (.A(_09423_),
    .ZN(_09806_));
 OAI21_X1 _19466_ (.A(_08565_),
    .B1(_08697_),
    .B2(_08606_),
    .ZN(_09807_));
 NAND2_X1 _19467_ (.A1(_08565_),
    .A2(_08718_),
    .ZN(_09808_));
 AND4_X1 _19468_ (.A1(_09806_),
    .A2(_09807_),
    .A3(_09553_),
    .A4(_09808_),
    .ZN(_09809_));
 AND2_X1 _19469_ (.A1(_08631_),
    .A2(_08651_),
    .ZN(_09810_));
 OAI21_X1 _19470_ (.A(_08549_),
    .B1(_08698_),
    .B2(_09810_),
    .ZN(_09811_));
 NAND3_X1 _19471_ (.A1(_08588_),
    .A2(_08549_),
    .A3(_08590_),
    .ZN(_09812_));
 AND4_X1 _19472_ (.A1(_08554_),
    .A2(_09809_),
    .A3(_09811_),
    .A4(_09812_),
    .ZN(_09813_));
 AOI21_X1 _19473_ (.A(_08560_),
    .B1(_09599_),
    .B2(_08680_),
    .ZN(_09814_));
 AOI21_X1 _19474_ (.A(_08560_),
    .B1(_08528_),
    .B2(_09585_),
    .ZN(_09815_));
 NOR3_X1 _19475_ (.A1(_09814_),
    .A2(_09815_),
    .A3(_09413_),
    .ZN(_09816_));
 OAI21_X1 _19476_ (.A(_08664_),
    .B1(_08708_),
    .B2(_08578_),
    .ZN(_09817_));
 OAI21_X1 _19477_ (.A(_08663_),
    .B1(_08797_),
    .B2(_08607_),
    .ZN(_09818_));
 OAI21_X1 _19478_ (.A(_08664_),
    .B1(_08544_),
    .B2(_08553_),
    .ZN(_09819_));
 AND4_X1 _19479_ (.A1(_09816_),
    .A2(_09817_),
    .A3(_09818_),
    .A4(_09819_),
    .ZN(_09820_));
 NAND3_X1 _19480_ (.A1(_08599_),
    .A2(_08526_),
    .A3(_08614_),
    .ZN(_09821_));
 NAND4_X1 _19481_ (.A1(_08657_),
    .A2(_08633_),
    .A3(_08593_),
    .A4(_08579_),
    .ZN(_09822_));
 AND3_X1 _19482_ (.A1(_09821_),
    .A2(_09397_),
    .A3(_09822_),
    .ZN(_09823_));
 OAI21_X1 _19483_ (.A(_08542_),
    .B1(_08536_),
    .B2(_08640_),
    .ZN(_09824_));
 NAND2_X1 _19484_ (.A1(_08640_),
    .A2(_08599_),
    .ZN(_09825_));
 NAND4_X1 _19485_ (.A1(_08631_),
    .A2(_08540_),
    .A3(_08509_),
    .A4(_08633_),
    .ZN(_09826_));
 AND3_X1 _19486_ (.A1(_08799_),
    .A2(_09825_),
    .A3(_09826_),
    .ZN(_09827_));
 OAI21_X1 _19487_ (.A(_08542_),
    .B1(_08685_),
    .B2(_08611_),
    .ZN(_09828_));
 AND4_X1 _19488_ (.A1(_09823_),
    .A2(_09824_),
    .A3(_09827_),
    .A4(_09828_),
    .ZN(_09829_));
 NAND2_X1 _19489_ (.A1(_08586_),
    .A2(_08698_),
    .ZN(_09830_));
 OAI21_X1 _19490_ (.A(_08585_),
    .B1(_08689_),
    .B2(_08544_),
    .ZN(_09831_));
 NAND3_X1 _19491_ (.A1(_08670_),
    .A2(_08731_),
    .A3(_08636_),
    .ZN(_09832_));
 NAND2_X1 _19492_ (.A1(_08636_),
    .A2(_08640_),
    .ZN(_09833_));
 AND4_X1 _19493_ (.A1(_09830_),
    .A2(_09831_),
    .A3(_09832_),
    .A4(_09833_),
    .ZN(_09834_));
 NAND4_X1 _19494_ (.A1(_09813_),
    .A2(_09820_),
    .A3(_09829_),
    .A4(_09834_),
    .ZN(_09835_));
 NOR2_X2 _19495_ (.A1(_09805_),
    .A2(_09835_),
    .ZN(_09836_));
 AND2_X1 _19496_ (.A1(_07117_),
    .A2(_06853_),
    .ZN(_09837_));
 INV_X1 _19497_ (.A(_09837_),
    .ZN(_09838_));
 AOI21_X1 _19498_ (.A(_07685_),
    .B1(_09314_),
    .B2(_09838_),
    .ZN(_09839_));
 AOI211_X1 _19499_ (.A(_09515_),
    .B(_09839_),
    .C1(_08422_),
    .C2(_08337_),
    .ZN(_09840_));
 AND2_X1 _19500_ (.A1(_07073_),
    .A2(_09313_),
    .ZN(_09841_));
 AND2_X1 _19501_ (.A1(_08091_),
    .A2(_16714_),
    .ZN(_09842_));
 AND2_X1 _19502_ (.A1(_07073_),
    .A2(_09842_),
    .ZN(_09843_));
 AOI221_X4 _19503_ (.A(_09841_),
    .B1(_09263_),
    .B2(_07084_),
    .C1(_06908_),
    .C2(_09843_),
    .ZN(_09844_));
 AND4_X1 _19504_ (.A1(_09334_),
    .A2(_09840_),
    .A3(_09506_),
    .A4(_09844_),
    .ZN(_09845_));
 NAND2_X1 _19505_ (.A1(_07348_),
    .A2(_06732_),
    .ZN(_09846_));
 NAND4_X1 _19506_ (.A1(_08069_),
    .A2(_07598_),
    .A3(_08113_),
    .A4(_08463_),
    .ZN(_09847_));
 OAI211_X1 _19507_ (.A(_09846_),
    .B(_09847_),
    .C1(_08482_),
    .C2(_07488_),
    .ZN(_09848_));
 AOI21_X1 _19508_ (.A(_07488_),
    .B1(_08318_),
    .B2(_08327_),
    .ZN(_09849_));
 AND4_X1 _19509_ (.A1(_08102_),
    .A2(_08478_),
    .A3(_08113_),
    .A4(_08463_),
    .ZN(_09850_));
 NOR3_X1 _19510_ (.A1(_09848_),
    .A2(_09849_),
    .A3(_09850_),
    .ZN(_09851_));
 OAI21_X1 _19511_ (.A(_08025_),
    .B1(_07981_),
    .B2(_07348_),
    .ZN(_09852_));
 NAND2_X1 _19512_ (.A1(_08025_),
    .A2(_06952_),
    .ZN(_09853_));
 OAI21_X1 _19513_ (.A(_08014_),
    .B1(_07029_),
    .B2(_06776_),
    .ZN(_09854_));
 AND3_X1 _19514_ (.A1(_09852_),
    .A2(_09853_),
    .A3(_09854_),
    .ZN(_09855_));
 AND2_X1 _19515_ (.A1(_09313_),
    .A2(_07828_),
    .ZN(_09856_));
 AND2_X1 _19516_ (.A1(_07532_),
    .A2(_07828_),
    .ZN(_09857_));
 AOI211_X1 _19517_ (.A(_09856_),
    .B(_09857_),
    .C1(_08498_),
    .C2(_07839_),
    .ZN(_09858_));
 NAND3_X1 _19518_ (.A1(_07444_),
    .A2(_09325_),
    .A3(_07400_),
    .ZN(_09859_));
 NAND2_X1 _19519_ (.A1(_07348_),
    .A2(_07400_),
    .ZN(_09860_));
 AND2_X1 _19520_ (.A1(_09859_),
    .A2(_09860_),
    .ZN(_09861_));
 AND4_X1 _19521_ (.A1(_09851_),
    .A2(_09855_),
    .A3(_09858_),
    .A4(_09861_),
    .ZN(_09862_));
 AOI211_X1 _19522_ (.A(_06842_),
    .B(_09311_),
    .C1(_08459_),
    .C2(_08102_),
    .ZN(_09863_));
 AND4_X1 _19523_ (.A1(_07161_),
    .A2(_08080_),
    .A3(_08233_),
    .A4(_08113_),
    .ZN(_09864_));
 AND4_X1 _19524_ (.A1(_06875_),
    .A2(_08461_),
    .A3(_08080_),
    .A4(_08113_),
    .ZN(_09865_));
 NOR4_X1 _19525_ (.A1(_09863_),
    .A2(_09312_),
    .A3(_09864_),
    .A4(_09865_),
    .ZN(_09866_));
 INV_X1 _19526_ (.A(_09331_),
    .ZN(_09867_));
 NAND2_X1 _19527_ (.A1(_08156_),
    .A2(_08233_),
    .ZN(_09868_));
 NAND2_X1 _19528_ (.A1(_08156_),
    .A2(_09289_),
    .ZN(_09869_));
 OAI21_X1 _19529_ (.A(_08156_),
    .B1(_08498_),
    .B2(_08451_),
    .ZN(_09870_));
 AND4_X1 _19530_ (.A1(_09867_),
    .A2(_09868_),
    .A3(_09869_),
    .A4(_09870_),
    .ZN(_09871_));
 NAND4_X1 _19531_ (.A1(_09845_),
    .A2(_09862_),
    .A3(_09866_),
    .A4(_09871_),
    .ZN(_09872_));
 INV_X1 _19532_ (.A(_09356_),
    .ZN(_09873_));
 AOI21_X1 _19533_ (.A(_09346_),
    .B1(_08468_),
    .B2(_09287_),
    .ZN(_09874_));
 AND4_X1 _19534_ (.A1(_07194_),
    .A2(_08211_),
    .A3(_08403_),
    .A4(_08113_),
    .ZN(_09875_));
 NOR3_X1 _19535_ (.A1(_09874_),
    .A2(_09462_),
    .A3(_09875_),
    .ZN(_09876_));
 AND2_X1 _19536_ (.A1(_09348_),
    .A2(_09352_),
    .ZN(_09877_));
 INV_X1 _19537_ (.A(_09877_),
    .ZN(_09878_));
 OAI211_X1 _19538_ (.A(_08200_),
    .B(_08222_),
    .C1(_08498_),
    .C2(_06776_),
    .ZN(_09879_));
 AND4_X1 _19539_ (.A1(_09873_),
    .A2(_09876_),
    .A3(_09878_),
    .A4(_09879_),
    .ZN(_09880_));
 AND4_X1 _19540_ (.A1(_07183_),
    .A2(_08211_),
    .A3(_08403_),
    .A4(_07554_),
    .ZN(_09881_));
 AND4_X1 _19541_ (.A1(_06754_),
    .A2(_08211_),
    .A3(_07183_),
    .A4(_07554_),
    .ZN(_09882_));
 AOI211_X1 _19542_ (.A(_09881_),
    .B(_09882_),
    .C1(_07315_),
    .C2(_09272_),
    .ZN(_09883_));
 AND3_X1 _19543_ (.A1(_09313_),
    .A2(_08211_),
    .A3(_07554_),
    .ZN(_09884_));
 AND3_X1 _19544_ (.A1(_09359_),
    .A2(_09325_),
    .A3(_07315_),
    .ZN(_09885_));
 AOI211_X1 _19545_ (.A(_09884_),
    .B(_09885_),
    .C1(_09456_),
    .C2(_07315_),
    .ZN(_09886_));
 NAND2_X1 _19546_ (.A1(_09322_),
    .A2(_07663_),
    .ZN(_09887_));
 OAI21_X1 _19547_ (.A(_08485_),
    .B1(_09887_),
    .B2(_06776_),
    .ZN(_09888_));
 OAI21_X1 _19548_ (.A(_08485_),
    .B1(_09327_),
    .B2(_07609_),
    .ZN(_09889_));
 AND4_X1 _19549_ (.A1(_09883_),
    .A2(_09886_),
    .A3(_09888_),
    .A4(_09889_),
    .ZN(_09890_));
 AOI211_X1 _19550_ (.A(_06842_),
    .B(_09261_),
    .C1(_08459_),
    .C2(_08102_),
    .ZN(_09891_));
 NAND2_X1 _19551_ (.A1(_07216_),
    .A2(_07565_),
    .ZN(_09892_));
 NAND3_X1 _19552_ (.A1(_07576_),
    .A2(_07150_),
    .A3(_07356_),
    .ZN(_09893_));
 OAI211_X1 _19553_ (.A(_09892_),
    .B(_09893_),
    .C1(_09287_),
    .C2(_09261_),
    .ZN(_09894_));
 OAI21_X1 _19554_ (.A(_08472_),
    .B1(_09322_),
    .B2(_09261_),
    .ZN(_09895_));
 NOR3_X1 _19555_ (.A1(_09891_),
    .A2(_09894_),
    .A3(_09895_),
    .ZN(_09896_));
 AND2_X1 _19556_ (.A1(_07784_),
    .A2(_07007_),
    .ZN(_09897_));
 AND2_X1 _19557_ (.A1(_07762_),
    .A2(_07007_),
    .ZN(_09898_));
 AND2_X1 _19558_ (.A1(_07532_),
    .A2(_07007_),
    .ZN(_09899_));
 NOR4_X1 _19559_ (.A1(_07018_),
    .A2(_09897_),
    .A3(_09898_),
    .A4(_09899_),
    .ZN(_09900_));
 OAI211_X1 _19560_ (.A(_08450_),
    .B(_08461_),
    .C1(_08459_),
    .C2(_08102_),
    .ZN(_09901_));
 OAI21_X1 _19561_ (.A(_08450_),
    .B1(_07348_),
    .B2(_09456_),
    .ZN(_09902_));
 AND4_X1 _19562_ (.A1(_09896_),
    .A2(_09900_),
    .A3(_09901_),
    .A4(_09902_),
    .ZN(_09903_));
 OAI21_X1 _19563_ (.A(_08491_),
    .B1(_09887_),
    .B2(_07532_),
    .ZN(_09904_));
 NAND2_X1 _19564_ (.A1(_07249_),
    .A2(_07378_),
    .ZN(_09905_));
 NAND2_X1 _19565_ (.A1(_09330_),
    .A2(_07227_),
    .ZN(_09906_));
 AND4_X1 _19566_ (.A1(_09281_),
    .A2(_09905_),
    .A3(_09284_),
    .A4(_09906_),
    .ZN(_09907_));
 AND4_X1 _19567_ (.A1(_07543_),
    .A2(_07183_),
    .A3(_08403_),
    .A4(_06699_),
    .ZN(_09908_));
 AND2_X1 _19568_ (.A1(_07238_),
    .A2(_08451_),
    .ZN(_09909_));
 AOI211_X1 _19569_ (.A(_09908_),
    .B(_09909_),
    .C1(_07249_),
    .C2(_07904_),
    .ZN(_09910_));
 OAI21_X1 _19570_ (.A(_08491_),
    .B1(_07948_),
    .B2(_09456_),
    .ZN(_09911_));
 AND4_X1 _19571_ (.A1(_09904_),
    .A2(_09907_),
    .A3(_09910_),
    .A4(_09911_),
    .ZN(_09912_));
 NAND4_X1 _19572_ (.A1(_09880_),
    .A2(_09890_),
    .A3(_09903_),
    .A4(_09912_),
    .ZN(_09913_));
 NOR2_X2 _19573_ (.A1(_09872_),
    .A2(_09913_),
    .ZN(_09914_));
 XOR2_X1 _19574_ (.A(_09836_),
    .B(_09914_),
    .Z(_09915_));
 NAND2_X1 _19575_ (.A1(_09116_),
    .A2(_08868_),
    .ZN(_09916_));
 NOR2_X1 _19576_ (.A1(_08866_),
    .A2(_09916_),
    .ZN(_09917_));
 AOI211_X1 _19577_ (.A(_08880_),
    .B(_09917_),
    .C1(_08998_),
    .C2(_09075_),
    .ZN(_09918_));
 AND4_X1 _19578_ (.A1(_08825_),
    .A2(_08864_),
    .A3(_08874_),
    .A4(_09115_),
    .ZN(_09919_));
 AND4_X1 _19579_ (.A1(_08825_),
    .A2(_08913_),
    .A3(_08858_),
    .A4(_08842_),
    .ZN(_09920_));
 AOI211_X1 _19580_ (.A(_09919_),
    .B(_09920_),
    .C1(_08904_),
    .C2(_09075_),
    .ZN(_09921_));
 OAI21_X1 _19581_ (.A(_08888_),
    .B1(_09074_),
    .B2(_08989_),
    .ZN(_09922_));
 OAI21_X1 _19582_ (.A(_08888_),
    .B1(_09046_),
    .B2(_08945_),
    .ZN(_09923_));
 AND4_X1 _19583_ (.A1(_09918_),
    .A2(_09921_),
    .A3(_09922_),
    .A4(_09923_),
    .ZN(_09924_));
 NOR2_X1 _19584_ (.A1(_08984_),
    .A2(_09115_),
    .ZN(_09925_));
 OAI21_X1 _19585_ (.A(_09106_),
    .B1(_09925_),
    .B2(_09095_),
    .ZN(_09926_));
 NAND2_X1 _19586_ (.A1(_09106_),
    .A2(_08943_),
    .ZN(_09927_));
 NAND2_X1 _19587_ (.A1(_08906_),
    .A2(_08986_),
    .ZN(_09928_));
 AND3_X1 _19588_ (.A1(_08912_),
    .A2(_09927_),
    .A3(_09928_),
    .ZN(_09929_));
 OAI21_X1 _19589_ (.A(_09720_),
    .B1(_08882_),
    .B2(_08904_),
    .ZN(_09930_));
 OAI21_X1 _19590_ (.A(_09720_),
    .B1(_09077_),
    .B2(_09710_),
    .ZN(_09931_));
 AND4_X1 _19591_ (.A1(_09926_),
    .A2(_09929_),
    .A3(_09930_),
    .A4(_09931_),
    .ZN(_09932_));
 OAI21_X1 _19592_ (.A(_08941_),
    .B1(_08986_),
    .B2(_08838_),
    .ZN(_09933_));
 OAI21_X1 _19593_ (.A(_08941_),
    .B1(_08903_),
    .B2(_08909_),
    .ZN(_09934_));
 OAI21_X1 _19594_ (.A(_08936_),
    .B1(_08986_),
    .B2(_09710_),
    .ZN(_09935_));
 OAI21_X1 _19595_ (.A(_08936_),
    .B1(_08903_),
    .B2(_08945_),
    .ZN(_09936_));
 AND4_X1 _19596_ (.A1(_09933_),
    .A2(_09934_),
    .A3(_09935_),
    .A4(_09936_),
    .ZN(_09937_));
 INV_X1 _19597_ (.A(_09059_),
    .ZN(_09938_));
 INV_X1 _19598_ (.A(_09070_),
    .ZN(_09939_));
 OAI21_X1 _19599_ (.A(_08834_),
    .B1(_08954_),
    .B2(_09014_),
    .ZN(_09940_));
 AND4_X1 _19600_ (.A1(_08851_),
    .A2(_09939_),
    .A3(_08856_),
    .A4(_09940_),
    .ZN(_09941_));
 NAND2_X1 _19601_ (.A1(_09730_),
    .A2(_09116_),
    .ZN(_09942_));
 NAND3_X1 _19602_ (.A1(_08829_),
    .A2(_09029_),
    .A3(_09115_),
    .ZN(_09943_));
 AND2_X1 _19603_ (.A1(_09942_),
    .A2(_09943_),
    .ZN(_09944_));
 NAND3_X1 _19604_ (.A1(_09122_),
    .A2(_08867_),
    .A3(_08829_),
    .ZN(_09945_));
 AND4_X1 _19605_ (.A1(_09938_),
    .A2(_09941_),
    .A3(_09944_),
    .A4(_09945_),
    .ZN(_09946_));
 NAND4_X1 _19606_ (.A1(_09924_),
    .A2(_09932_),
    .A3(_09937_),
    .A4(_09946_),
    .ZN(_09947_));
 OAI21_X1 _19607_ (.A(_09087_),
    .B1(_08903_),
    .B2(_08969_),
    .ZN(_09948_));
 AND2_X1 _19608_ (.A1(_08938_),
    .A2(_08982_),
    .ZN(_09949_));
 AND2_X1 _19609_ (.A1(_08982_),
    .A2(_08987_),
    .ZN(_09950_));
 AND2_X1 _19610_ (.A1(_08976_),
    .A2(_08945_),
    .ZN(_09951_));
 NOR4_X1 _19611_ (.A1(_09949_),
    .A2(_09950_),
    .A3(_09951_),
    .A4(_08978_),
    .ZN(_09952_));
 NAND4_X1 _19612_ (.A1(_08886_),
    .A2(_08843_),
    .A3(_08950_),
    .A4(_08973_),
    .ZN(_09953_));
 OAI21_X1 _19613_ (.A(_09087_),
    .B1(_09017_),
    .B2(_08998_),
    .ZN(_09954_));
 AND4_X1 _19614_ (.A1(_09948_),
    .A2(_09952_),
    .A3(_09953_),
    .A4(_09954_),
    .ZN(_09955_));
 OR2_X1 _19615_ (.A1(_09109_),
    .A2(_09916_),
    .ZN(_09956_));
 AND2_X1 _19616_ (.A1(_09007_),
    .A2(_08855_),
    .ZN(_09957_));
 AND2_X1 _19617_ (.A1(_09007_),
    .A2(_08850_),
    .ZN(_09958_));
 AND2_X1 _19618_ (.A1(_09007_),
    .A2(_08915_),
    .ZN(_09959_));
 AND2_X1 _19619_ (.A1(_09007_),
    .A2(_08969_),
    .ZN(_09960_));
 NOR4_X1 _19620_ (.A1(_09957_),
    .A2(_09958_),
    .A3(_09959_),
    .A4(_09960_),
    .ZN(_09961_));
 OAI21_X1 _19621_ (.A(_09005_),
    .B1(_08998_),
    .B2(_08987_),
    .ZN(_09962_));
 OAI211_X1 _19622_ (.A(_09005_),
    .B(_16794_),
    .C1(_08845_),
    .C2(_08816_),
    .ZN(_09963_));
 AND4_X1 _19623_ (.A1(_09956_),
    .A2(_09961_),
    .A3(_09962_),
    .A4(_09963_),
    .ZN(_09964_));
 OAI211_X1 _19624_ (.A(_09053_),
    .B(_09029_),
    .C1(_08973_),
    .C2(_08878_),
    .ZN(_09965_));
 NAND2_X1 _19625_ (.A1(_08959_),
    .A2(_09965_),
    .ZN(_09966_));
 OAI211_X1 _19626_ (.A(_08972_),
    .B(_09029_),
    .C1(_08823_),
    .C2(_09115_),
    .ZN(_09967_));
 OAI21_X1 _19627_ (.A(_08972_),
    .B1(_08943_),
    .B2(_08915_),
    .ZN(_09968_));
 OAI21_X1 _19628_ (.A(_08952_),
    .B1(_09009_),
    .B2(_08909_),
    .ZN(_09969_));
 NAND4_X1 _19629_ (.A1(_09967_),
    .A2(_09968_),
    .A3(_09969_),
    .A4(_09696_),
    .ZN(_09970_));
 AND2_X1 _19630_ (.A1(_09053_),
    .A2(_08915_),
    .ZN(_09971_));
 NOR4_X1 _19631_ (.A1(_09966_),
    .A2(_09970_),
    .A3(_08963_),
    .A4(_09971_),
    .ZN(_09972_));
 OAI21_X1 _19632_ (.A(_09026_),
    .B1(_09095_),
    .B2(_08903_),
    .ZN(_09973_));
 NAND3_X1 _19633_ (.A1(_08933_),
    .A2(_09003_),
    .A3(_08864_),
    .ZN(_09974_));
 NAND2_X1 _19634_ (.A1(_09026_),
    .A2(_08911_),
    .ZN(_09975_));
 AND4_X1 _19635_ (.A1(_09723_),
    .A2(_09973_),
    .A3(_09974_),
    .A4(_09975_),
    .ZN(_09976_));
 AND2_X1 _19636_ (.A1(_08850_),
    .A2(_09020_),
    .ZN(_09977_));
 AND2_X1 _19637_ (.A1(_09020_),
    .A2(_09009_),
    .ZN(_09978_));
 AND4_X1 _19638_ (.A1(_08886_),
    .A2(_08874_),
    .A3(_09115_),
    .A4(_09003_),
    .ZN(_09979_));
 NOR4_X1 _19639_ (.A1(_09022_),
    .A2(_09977_),
    .A3(_09978_),
    .A4(_09979_),
    .ZN(_09980_));
 OAI211_X1 _19640_ (.A(_09031_),
    .B(_09107_),
    .C1(_08844_),
    .C2(_08845_),
    .ZN(_09981_));
 AND4_X1 _19641_ (.A1(_09100_),
    .A2(_09976_),
    .A3(_09980_),
    .A4(_09981_),
    .ZN(_09982_));
 NAND4_X1 _19642_ (.A1(_09955_),
    .A2(_09964_),
    .A3(_09972_),
    .A4(_09982_),
    .ZN(_09983_));
 NOR2_X2 _19643_ (.A1(_09947_),
    .A2(_09983_),
    .ZN(_09984_));
 XOR2_X1 _19644_ (.A(_09984_),
    .B(_09035_),
    .Z(_09985_));
 XNOR2_X1 _19645_ (.A(_09915_),
    .B(_09985_),
    .ZN(_09986_));
 XNOR2_X1 _19646_ (.A(_09603_),
    .B(_08811_),
    .ZN(_09987_));
 NAND2_X1 _19647_ (.A1(_06171_),
    .A2(_06490_),
    .ZN(_09988_));
 NAND4_X1 _19648_ (.A1(_05687_),
    .A2(_04439_),
    .A3(_04735_),
    .A4(_06149_),
    .ZN(_09989_));
 AND2_X1 _19649_ (.A1(_06204_),
    .A2(_09989_),
    .ZN(_09990_));
 NAND2_X1 _19650_ (.A1(_06171_),
    .A2(_04307_),
    .ZN(_09991_));
 NAND4_X1 _19651_ (.A1(_06193_),
    .A2(_09988_),
    .A3(_09990_),
    .A4(_09991_),
    .ZN(_09992_));
 AND4_X1 _19652_ (.A1(_06325_),
    .A2(_04950_),
    .A3(_06149_),
    .A4(_04592_),
    .ZN(_09993_));
 OR2_X1 _19653_ (.A1(_09211_),
    .A2(_09213_),
    .ZN(_09994_));
 NAND2_X1 _19654_ (.A1(_04395_),
    .A2(_06270_),
    .ZN(_09995_));
 NAND2_X1 _19655_ (.A1(_04636_),
    .A2(_06270_),
    .ZN(_09996_));
 INV_X1 _19656_ (.A(_06281_),
    .ZN(_09997_));
 OAI221_X1 _19657_ (.A(_09995_),
    .B1(_09996_),
    .B2(_06325_),
    .C1(_09997_),
    .C2(_06105_),
    .ZN(_09998_));
 NOR4_X1 _19658_ (.A1(_09992_),
    .A2(_09993_),
    .A3(_09994_),
    .A4(_09998_),
    .ZN(_09999_));
 OAI211_X1 _19659_ (.A(_04461_),
    .B(_09158_),
    .C1(_04395_),
    .C2(_05096_),
    .ZN(_10000_));
 INV_X1 _19660_ (.A(_04636_),
    .ZN(_10001_));
 OAI21_X1 _19661_ (.A(_10000_),
    .B1(_10001_),
    .B2(_09197_),
    .ZN(_10002_));
 INV_X1 _19662_ (.A(_04855_),
    .ZN(_10003_));
 AOI21_X1 _19663_ (.A(_09197_),
    .B1(_05918_),
    .B2(_10003_),
    .ZN(_10004_));
 AND2_X1 _19664_ (.A1(_05045_),
    .A2(_09182_),
    .ZN(_10005_));
 NOR4_X1 _19665_ (.A1(_10002_),
    .A2(_10004_),
    .A3(_09203_),
    .A4(_10005_),
    .ZN(_10006_));
 OAI211_X1 _19666_ (.A(_04614_),
    .B(_04950_),
    .C1(_06314_),
    .C2(_05203_),
    .ZN(_10007_));
 AND2_X1 _19667_ (.A1(_04384_),
    .A2(_05116_),
    .ZN(_10008_));
 OAI21_X1 _19668_ (.A(_04614_),
    .B1(_09615_),
    .B2(_10008_),
    .ZN(_10009_));
 AND4_X1 _19669_ (.A1(_09188_),
    .A2(_10006_),
    .A3(_10007_),
    .A4(_10009_),
    .ZN(_10010_));
 AND2_X1 _19670_ (.A1(_04669_),
    .A2(_05116_),
    .ZN(_10011_));
 OAI21_X1 _19671_ (.A(_04888_),
    .B1(_09623_),
    .B2(_10011_),
    .ZN(_10012_));
 OAI211_X1 _19672_ (.A(_10012_),
    .B(_09659_),
    .C1(_06248_),
    .C2(_09193_),
    .ZN(_10013_));
 AND2_X1 _19673_ (.A1(_04494_),
    .A2(_09178_),
    .ZN(_10014_));
 OAI21_X1 _19674_ (.A(_04494_),
    .B1(_09623_),
    .B2(_05159_),
    .ZN(_10015_));
 NAND2_X1 _19675_ (.A1(_04494_),
    .A2(_05082_),
    .ZN(_10016_));
 NAND2_X1 _19676_ (.A1(_10015_),
    .A2(_10016_),
    .ZN(_10017_));
 NOR4_X1 _19677_ (.A1(_10013_),
    .A2(_09206_),
    .A3(_10014_),
    .A4(_10017_),
    .ZN(_10018_));
 NAND2_X1 _19678_ (.A1(_06446_),
    .A2(_09623_),
    .ZN(_10019_));
 OAI21_X1 _19679_ (.A(_06567_),
    .B1(_04340_),
    .B2(_04746_),
    .ZN(_10020_));
 OAI21_X1 _19680_ (.A(_06446_),
    .B1(_05120_),
    .B2(_04855_),
    .ZN(_10021_));
 NAND2_X1 _19681_ (.A1(_06490_),
    .A2(_06567_),
    .ZN(_10022_));
 AND4_X1 _19682_ (.A1(_10019_),
    .A2(_10020_),
    .A3(_10021_),
    .A4(_10022_),
    .ZN(_10023_));
 NAND4_X1 _19683_ (.A1(_09999_),
    .A2(_10010_),
    .A3(_10018_),
    .A4(_10023_),
    .ZN(_10024_));
 NAND4_X1 _19684_ (.A1(_05324_),
    .A2(_06325_),
    .A3(_04833_),
    .A4(_04950_),
    .ZN(_10025_));
 NAND2_X1 _19685_ (.A1(_05291_),
    .A2(_05096_),
    .ZN(_10026_));
 NOR2_X1 _19686_ (.A1(_05269_),
    .A2(_09642_),
    .ZN(_10027_));
 AND2_X1 _19687_ (.A1(_05599_),
    .A2(_05258_),
    .ZN(_10028_));
 INV_X1 _19688_ (.A(_10028_),
    .ZN(_10029_));
 AND4_X1 _19689_ (.A1(_10026_),
    .A2(_10027_),
    .A3(_09177_),
    .A4(_10029_),
    .ZN(_10030_));
 OAI211_X1 _19690_ (.A(_05401_),
    .B(_06303_),
    .C1(_06314_),
    .C2(_05203_),
    .ZN(_10031_));
 AND4_X1 _19691_ (.A1(_05137_),
    .A2(_05324_),
    .A3(_05797_),
    .A4(_04833_),
    .ZN(_10032_));
 AOI211_X1 _19692_ (.A(_10032_),
    .B(_09150_),
    .C1(_05401_),
    .C2(_06138_),
    .ZN(_10033_));
 AND4_X1 _19693_ (.A1(_10025_),
    .A2(_10030_),
    .A3(_10031_),
    .A4(_10033_),
    .ZN(_10034_));
 OAI211_X1 _19694_ (.A(_09251_),
    .B(_05863_),
    .C1(_04959_),
    .C2(_06325_),
    .ZN(_10035_));
 OAI21_X1 _19695_ (.A(_09251_),
    .B1(_04263_),
    .B2(_04307_),
    .ZN(_10036_));
 OAI211_X1 _19696_ (.A(_09251_),
    .B(_04950_),
    .C1(_05368_),
    .C2(_05313_),
    .ZN(_10037_));
 OAI21_X1 _19697_ (.A(_09251_),
    .B1(_06490_),
    .B2(_05159_),
    .ZN(_10038_));
 NAND4_X1 _19698_ (.A1(_10035_),
    .A2(_10036_),
    .A3(_10037_),
    .A4(_10038_),
    .ZN(_10039_));
 OAI211_X1 _19699_ (.A(_09246_),
    .B(_05863_),
    .C1(_06314_),
    .C2(_06325_),
    .ZN(_10040_));
 OAI21_X1 _19700_ (.A(_10040_),
    .B1(_09186_),
    .B2(_09248_),
    .ZN(_10041_));
 OAI21_X1 _19701_ (.A(_06050_),
    .B1(_09248_),
    .B2(_05456_),
    .ZN(_10042_));
 AOI21_X1 _19702_ (.A(_09248_),
    .B1(_09198_),
    .B2(_09194_),
    .ZN(_10043_));
 NOR4_X1 _19703_ (.A1(_10039_),
    .A2(_10041_),
    .A3(_10042_),
    .A4(_10043_),
    .ZN(_10044_));
 NAND2_X1 _19704_ (.A1(_09198_),
    .A2(_09194_),
    .ZN(_10045_));
 OAI21_X1 _19705_ (.A(_05632_),
    .B1(_10045_),
    .B2(_05120_),
    .ZN(_10046_));
 NAND3_X1 _19706_ (.A1(_10046_),
    .A2(_05643_),
    .A3(_09618_),
    .ZN(_10047_));
 OAI21_X1 _19707_ (.A(_05786_),
    .B1(_05017_),
    .B2(_04778_),
    .ZN(_10048_));
 NAND2_X1 _19708_ (.A1(_04746_),
    .A2(_05786_),
    .ZN(_10049_));
 NAND2_X1 _19709_ (.A1(_10048_),
    .A2(_10049_),
    .ZN(_10050_));
 AOI21_X1 _19710_ (.A(_09238_),
    .B1(_10001_),
    .B2(_05170_),
    .ZN(_10051_));
 AOI21_X1 _19711_ (.A(_09238_),
    .B1(_06105_),
    .B2(_04526_),
    .ZN(_10052_));
 NOR4_X1 _19712_ (.A1(_10047_),
    .A2(_10050_),
    .A3(_10051_),
    .A4(_10052_),
    .ZN(_10053_));
 OAI21_X1 _19713_ (.A(_05522_),
    .B1(_09639_),
    .B2(_09182_),
    .ZN(_10054_));
 OAI211_X1 _19714_ (.A(_10054_),
    .B(_09632_),
    .C1(_09194_),
    .C2(_09168_),
    .ZN(_10055_));
 AND2_X1 _19715_ (.A1(_09169_),
    .A2(_05214_),
    .ZN(_10056_));
 AOI21_X1 _19716_ (.A(_05114_),
    .B1(_05434_),
    .B2(_10003_),
    .ZN(_10057_));
 NOR4_X1 _19717_ (.A1(_10055_),
    .A2(_10056_),
    .A3(_09160_),
    .A4(_10057_),
    .ZN(_10058_));
 NAND4_X1 _19718_ (.A1(_10034_),
    .A2(_10044_),
    .A3(_10053_),
    .A4(_10058_),
    .ZN(_10059_));
 NOR2_X2 _19719_ (.A1(_10024_),
    .A2(_10059_),
    .ZN(_10060_));
 XNOR2_X1 _19720_ (.A(_09987_),
    .B(_10060_),
    .ZN(_10061_));
 XNOR2_X1 _19721_ (.A(_09986_),
    .B(_10061_),
    .ZN(_10062_));
 XNOR2_X1 _19722_ (.A(_10062_),
    .B(_17092_),
    .ZN(_10063_));
 MUX2_X1 _19723_ (.A(_09763_),
    .B(_10063_),
    .S(_09040_),
    .Z(_00727_));
 XOR2_X1 _19724_ (.A(_17093_),
    .B(_17007_),
    .Z(_10064_));
 XNOR2_X1 _19725_ (.A(_09836_),
    .B(_08811_),
    .ZN(_10065_));
 AND2_X1 _19726_ (.A1(_05148_),
    .A2(_06545_),
    .ZN(_10066_));
 AND3_X1 _19727_ (.A1(_06556_),
    .A2(_05313_),
    .A3(_04669_),
    .ZN(_10067_));
 AOI211_X1 _19728_ (.A(_10066_),
    .B(_10067_),
    .C1(_06567_),
    .C2(_05379_),
    .ZN(_10068_));
 OAI21_X1 _19729_ (.A(_06446_),
    .B1(_06138_),
    .B2(_05797_),
    .ZN(_10069_));
 AND4_X1 _19730_ (.A1(_06435_),
    .A2(_10068_),
    .A3(_09221_),
    .A4(_10069_),
    .ZN(_10070_));
 AND2_X1 _19731_ (.A1(_06171_),
    .A2(_09615_),
    .ZN(_10071_));
 INV_X1 _19732_ (.A(_10071_),
    .ZN(_10072_));
 AND2_X1 _19733_ (.A1(_06171_),
    .A2(_05017_),
    .ZN(_10073_));
 INV_X1 _19734_ (.A(_10073_),
    .ZN(_10074_));
 NAND2_X1 _19735_ (.A1(_05379_),
    .A2(_06160_),
    .ZN(_10075_));
 OAI21_X1 _19736_ (.A(_06171_),
    .B1(_04395_),
    .B2(_06490_),
    .ZN(_10076_));
 NAND4_X1 _19737_ (.A1(_10072_),
    .A2(_10074_),
    .A3(_10075_),
    .A4(_10076_),
    .ZN(_10077_));
 NOR2_X1 _19738_ (.A1(_09997_),
    .A2(_06523_),
    .ZN(_10078_));
 AND3_X1 _19739_ (.A1(_06281_),
    .A2(_04735_),
    .A3(_04669_),
    .ZN(_10079_));
 OR2_X1 _19740_ (.A1(_09653_),
    .A2(_10079_),
    .ZN(_10080_));
 NOR4_X1 _19741_ (.A1(_10077_),
    .A2(_10078_),
    .A3(_10080_),
    .A4(_09212_),
    .ZN(_10081_));
 OAI21_X1 _19742_ (.A(_04494_),
    .B1(_05017_),
    .B2(_05445_),
    .ZN(_10082_));
 OAI211_X1 _19743_ (.A(_04494_),
    .B(_05797_),
    .C1(_04959_),
    .C2(_05203_),
    .ZN(_10083_));
 NAND4_X1 _19744_ (.A1(_04285_),
    .A2(_10016_),
    .A3(_10082_),
    .A4(_10083_),
    .ZN(_10084_));
 AOI21_X1 _19745_ (.A(_09193_),
    .B1(_10001_),
    .B2(_05170_),
    .ZN(_10085_));
 AND3_X1 _19746_ (.A1(_04844_),
    .A2(_04899_),
    .A3(_04669_),
    .ZN(_10086_));
 NAND2_X1 _19747_ (.A1(_04888_),
    .A2(_05064_),
    .ZN(_10087_));
 NAND2_X1 _19748_ (.A1(_04844_),
    .A2(_04307_),
    .ZN(_10088_));
 OAI211_X1 _19749_ (.A(_10087_),
    .B(_10088_),
    .C1(_09193_),
    .C2(_05456_),
    .ZN(_10089_));
 NOR4_X1 _19750_ (.A1(_10084_),
    .A2(_10085_),
    .A3(_10086_),
    .A4(_10089_),
    .ZN(_10090_));
 NAND3_X1 _19751_ (.A1(_05017_),
    .A2(_04592_),
    .A3(_04461_),
    .ZN(_10091_));
 OAI211_X1 _19752_ (.A(_04756_),
    .B(_10091_),
    .C1(_04800_),
    .C2(_09155_),
    .ZN(_10092_));
 NAND2_X1 _19753_ (.A1(_04997_),
    .A2(_09178_),
    .ZN(_10093_));
 NAND3_X1 _19754_ (.A1(_10093_),
    .A2(_05073_),
    .A3(_05103_),
    .ZN(_10094_));
 AOI21_X1 _19755_ (.A(_09197_),
    .B1(_09186_),
    .B2(_09183_),
    .ZN(_10095_));
 NOR4_X1 _19756_ (.A1(_10092_),
    .A2(_10094_),
    .A3(_10095_),
    .A4(_09184_),
    .ZN(_10096_));
 NAND4_X1 _19757_ (.A1(_10070_),
    .A2(_10081_),
    .A3(_10090_),
    .A4(_10096_),
    .ZN(_10097_));
 AND2_X1 _19758_ (.A1(_05302_),
    .A2(_05335_),
    .ZN(_10098_));
 NAND2_X1 _19759_ (.A1(_05291_),
    .A2(_05676_),
    .ZN(_10099_));
 AND3_X1 _19760_ (.A1(_09643_),
    .A2(_09176_),
    .A3(_10099_),
    .ZN(_10100_));
 OAI21_X1 _19761_ (.A(_05401_),
    .B1(_09178_),
    .B2(_05676_),
    .ZN(_10101_));
 OAI21_X1 _19762_ (.A(_05401_),
    .B1(_09169_),
    .B2(_09623_),
    .ZN(_10102_));
 AND4_X1 _19763_ (.A1(_10098_),
    .A2(_10100_),
    .A3(_10101_),
    .A4(_10102_),
    .ZN(_10103_));
 NAND4_X1 _19764_ (.A1(_05621_),
    .A2(_05643_),
    .A3(_09616_),
    .A4(_09618_),
    .ZN(_10104_));
 NAND2_X1 _19765_ (.A1(_09228_),
    .A2(_05786_),
    .ZN(_10105_));
 OAI21_X1 _19766_ (.A(_10105_),
    .B1(_09238_),
    .B2(_04789_),
    .ZN(_10106_));
 NAND3_X1 _19767_ (.A1(_05676_),
    .A2(_09158_),
    .A3(_05874_),
    .ZN(_10107_));
 OAI211_X1 _19768_ (.A(_10107_),
    .B(_09621_),
    .C1(_09155_),
    .C2(_05654_),
    .ZN(_10108_));
 NOR4_X1 _19769_ (.A1(_10104_),
    .A2(_09626_),
    .A3(_10106_),
    .A4(_10108_),
    .ZN(_10109_));
 OAI21_X1 _19770_ (.A(_09251_),
    .B1(_06534_),
    .B2(_04855_),
    .ZN(_10110_));
 OAI211_X1 _19771_ (.A(_09246_),
    .B(_16754_),
    .C1(_16753_),
    .C2(_05313_),
    .ZN(_10111_));
 OAI21_X1 _19772_ (.A(_09251_),
    .B1(_04537_),
    .B2(_05962_),
    .ZN(_10112_));
 AND4_X1 _19773_ (.A1(_06039_),
    .A2(_10110_),
    .A3(_10111_),
    .A4(_10112_),
    .ZN(_10113_));
 OAI21_X1 _19774_ (.A(_05522_),
    .B1(_04921_),
    .B2(_09182_),
    .ZN(_10114_));
 OAI21_X1 _19775_ (.A(_05214_),
    .B1(_04263_),
    .B2(_05017_),
    .ZN(_10115_));
 OAI21_X1 _19776_ (.A(_05214_),
    .B1(_09612_),
    .B2(_09182_),
    .ZN(_10116_));
 AND4_X1 _19777_ (.A1(_09166_),
    .A2(_10114_),
    .A3(_10115_),
    .A4(_10116_),
    .ZN(_10117_));
 NAND4_X1 _19778_ (.A1(_10103_),
    .A2(_10109_),
    .A3(_10113_),
    .A4(_10117_),
    .ZN(_10118_));
 NOR2_X2 _19779_ (.A1(_10097_),
    .A2(_10118_),
    .ZN(_10119_));
 XNOR2_X1 _19780_ (.A(_10065_),
    .B(_10119_),
    .ZN(_10120_));
 AND2_X1 _19781_ (.A1(_08564_),
    .A2(_08714_),
    .ZN(_10121_));
 INV_X1 _19782_ (.A(_10121_),
    .ZN(_10122_));
 NAND4_X1 _19783_ (.A1(_08665_),
    .A2(_08731_),
    .A3(_08632_),
    .A4(_08581_),
    .ZN(_10123_));
 OAI21_X1 _19784_ (.A(_08565_),
    .B1(_08568_),
    .B2(_08797_),
    .ZN(_10124_));
 AND4_X1 _19785_ (.A1(_09808_),
    .A2(_10122_),
    .A3(_10123_),
    .A4(_10124_),
    .ZN(_10125_));
 OAI21_X1 _19786_ (.A(_08549_),
    .B1(_08797_),
    .B2(_08607_),
    .ZN(_10126_));
 AND4_X1 _19787_ (.A1(_08653_),
    .A2(_08632_),
    .A3(_08593_),
    .A4(_08521_),
    .ZN(_10127_));
 AND2_X1 _19788_ (.A1(_08621_),
    .A2(_08548_),
    .ZN(_10128_));
 AOI211_X1 _19789_ (.A(_10127_),
    .B(_10128_),
    .C1(_08685_),
    .C2(_08549_),
    .ZN(_10129_));
 AND4_X1 _19790_ (.A1(_08766_),
    .A2(_10125_),
    .A3(_10126_),
    .A4(_10129_),
    .ZN(_10130_));
 OAI211_X1 _19791_ (.A(_08629_),
    .B(_08615_),
    .C1(_08618_),
    .C2(_08653_),
    .ZN(_10131_));
 OAI21_X1 _19792_ (.A(_10131_),
    .B1(_08678_),
    .B2(_08560_),
    .ZN(_10132_));
 NAND2_X1 _19793_ (.A1(_08704_),
    .A2(_08664_),
    .ZN(_10133_));
 NAND3_X1 _19794_ (.A1(_08724_),
    .A2(_08539_),
    .A3(_08632_),
    .ZN(_10134_));
 OAI211_X1 _19795_ (.A(_10133_),
    .B(_10134_),
    .C1(_09416_),
    .C2(_09581_),
    .ZN(_10135_));
 AOI21_X1 _19796_ (.A(_09416_),
    .B1(_08801_),
    .B2(_08694_),
    .ZN(_10136_));
 NOR4_X1 _19797_ (.A1(_10132_),
    .A2(_10135_),
    .A3(_10136_),
    .A4(_09411_),
    .ZN(_10137_));
 NAND2_X1 _19798_ (.A1(_08542_),
    .A2(_08553_),
    .ZN(_10138_));
 AND3_X1 _19799_ (.A1(_08640_),
    .A2(_08657_),
    .A3(_08539_),
    .ZN(_10139_));
 AOI211_X1 _19800_ (.A(_10139_),
    .B(_09399_),
    .C1(_08527_),
    .C2(_08542_),
    .ZN(_10140_));
 NAND2_X1 _19801_ (.A1(_09422_),
    .A2(_08599_),
    .ZN(_10141_));
 NAND2_X1 _19802_ (.A1(_08732_),
    .A2(_08622_),
    .ZN(_10142_));
 NAND2_X1 _19803_ (.A1(_08715_),
    .A2(_08622_),
    .ZN(_10143_));
 NAND3_X1 _19804_ (.A1(_08599_),
    .A2(_08653_),
    .A3(_08614_),
    .ZN(_10144_));
 AND4_X1 _19805_ (.A1(_10141_),
    .A2(_10142_),
    .A3(_10143_),
    .A4(_10144_),
    .ZN(_10145_));
 OAI211_X1 _19806_ (.A(_08542_),
    .B(_08615_),
    .C1(_09382_),
    .C2(_08574_),
    .ZN(_10146_));
 AND4_X1 _19807_ (.A1(_10138_),
    .A2(_10140_),
    .A3(_10145_),
    .A4(_10146_),
    .ZN(_10147_));
 NAND3_X1 _19808_ (.A1(_08586_),
    .A2(_08535_),
    .A3(_08531_),
    .ZN(_10148_));
 OAI211_X1 _19809_ (.A(_08625_),
    .B(_08614_),
    .C1(_08579_),
    .C2(_08574_),
    .ZN(_10149_));
 NAND4_X1 _19810_ (.A1(_08637_),
    .A2(_08642_),
    .A3(_08794_),
    .A4(_08657_),
    .ZN(_10150_));
 NAND4_X1 _19811_ (.A1(_08733_),
    .A2(_08526_),
    .A3(_08657_),
    .A4(_08642_),
    .ZN(_10151_));
 AND3_X1 _19812_ (.A1(_10149_),
    .A2(_10150_),
    .A3(_10151_),
    .ZN(_10152_));
 OAI21_X1 _19813_ (.A(_08586_),
    .B1(_09404_),
    .B2(_08672_),
    .ZN(_10153_));
 OAI211_X1 _19814_ (.A(_08657_),
    .B(_08581_),
    .C1(_08797_),
    .C2(_08607_),
    .ZN(_10154_));
 AND4_X1 _19815_ (.A1(_10148_),
    .A2(_10152_),
    .A3(_10153_),
    .A4(_10154_),
    .ZN(_10155_));
 NAND4_X1 _19816_ (.A1(_10130_),
    .A2(_10137_),
    .A3(_10147_),
    .A4(_10155_),
    .ZN(_10156_));
 OAI21_X1 _19817_ (.A(_08609_),
    .B1(_08705_),
    .B2(_08746_),
    .ZN(_10157_));
 OAI21_X1 _19818_ (.A(_08572_),
    .B1(_08594_),
    .B2(_08689_),
    .ZN(_10158_));
 AND4_X1 _19819_ (.A1(_08583_),
    .A2(_10157_),
    .A3(_09778_),
    .A4(_10158_),
    .ZN(_10159_));
 AND2_X1 _19820_ (.A1(_08519_),
    .A2(_08523_),
    .ZN(_10160_));
 INV_X1 _19821_ (.A(_10160_),
    .ZN(_10161_));
 OAI21_X1 _19822_ (.A(_08646_),
    .B1(_08797_),
    .B2(_08607_),
    .ZN(_10162_));
 OAI211_X1 _19823_ (.A(_10161_),
    .B(_10162_),
    .C1(_08528_),
    .C2(_08524_),
    .ZN(_10163_));
 AOI21_X1 _19824_ (.A(_08727_),
    .B1(_09796_),
    .B2(_09599_),
    .ZN(_10164_));
 AND4_X1 _19825_ (.A1(_09382_),
    .A2(_08581_),
    .A3(_08615_),
    .A4(_08675_),
    .ZN(_10165_));
 NAND2_X1 _19826_ (.A1(_08677_),
    .A2(_08682_),
    .ZN(_10166_));
 OAI21_X1 _19827_ (.A(_10166_),
    .B1(_08727_),
    .B2(_08802_),
    .ZN(_10167_));
 NOR4_X1 _19828_ (.A1(_10163_),
    .A2(_10164_),
    .A3(_10165_),
    .A4(_10167_),
    .ZN(_10168_));
 OAI211_X1 _19829_ (.A(_08703_),
    .B(_08733_),
    .C1(_09382_),
    .C2(_08794_),
    .ZN(_10169_));
 OAI21_X1 _19830_ (.A(_10169_),
    .B1(_09373_),
    .B2(_08768_),
    .ZN(_10170_));
 OAI211_X1 _19831_ (.A(_08741_),
    .B(_08742_),
    .C1(_09373_),
    .C2(_08557_),
    .ZN(_10171_));
 AOI21_X1 _19832_ (.A(_08529_),
    .B1(_09401_),
    .B2(_08557_),
    .ZN(_10172_));
 NOR4_X1 _19833_ (.A1(_10170_),
    .A2(_10171_),
    .A3(_09598_),
    .A4(_10172_),
    .ZN(_10173_));
 OAI21_X1 _19834_ (.A(_08650_),
    .B1(_08698_),
    .B2(_08606_),
    .ZN(_10174_));
 NAND2_X1 _19835_ (.A1(_08650_),
    .A2(_08708_),
    .ZN(_10175_));
 AND2_X1 _19836_ (.A1(_10174_),
    .A2(_10175_),
    .ZN(_10176_));
 OAI21_X1 _19837_ (.A(_08605_),
    .B1(_08714_),
    .B2(_08553_),
    .ZN(_10177_));
 OAI21_X1 _19838_ (.A(_08605_),
    .B1(_08732_),
    .B2(_08708_),
    .ZN(_10178_));
 AND4_X1 _19839_ (.A1(_09431_),
    .A2(_10176_),
    .A3(_10177_),
    .A4(_10178_),
    .ZN(_10179_));
 NAND4_X1 _19840_ (.A1(_10159_),
    .A2(_10168_),
    .A3(_10173_),
    .A4(_10179_),
    .ZN(_10180_));
 NOR2_X2 _19841_ (.A1(_10156_),
    .A2(_10180_),
    .ZN(_10181_));
 NAND2_X1 _19842_ (.A1(_08025_),
    .A2(_08451_),
    .ZN(_10182_));
 OAI21_X1 _19843_ (.A(_08014_),
    .B1(_09321_),
    .B2(_06952_),
    .ZN(_10183_));
 OAI21_X1 _19844_ (.A(_08014_),
    .B1(_08047_),
    .B2(_07348_),
    .ZN(_10184_));
 NAND3_X1 _19845_ (.A1(_07216_),
    .A2(_08189_),
    .A3(_08463_),
    .ZN(_10185_));
 AND4_X1 _19846_ (.A1(_10182_),
    .A2(_10183_),
    .A3(_10184_),
    .A4(_10185_),
    .ZN(_10186_));
 NAND2_X1 _19847_ (.A1(_07806_),
    .A2(_06732_),
    .ZN(_10187_));
 OAI21_X1 _19848_ (.A(_06732_),
    .B1(_07652_),
    .B2(_08473_),
    .ZN(_10188_));
 AND4_X1 _19849_ (.A1(_09522_),
    .A2(_10186_),
    .A3(_10187_),
    .A4(_10188_),
    .ZN(_10189_));
 OAI21_X1 _19850_ (.A(_07095_),
    .B1(_08047_),
    .B2(_07378_),
    .ZN(_10190_));
 NAND3_X1 _19851_ (.A1(_07084_),
    .A2(_08384_),
    .A3(_09325_),
    .ZN(_10191_));
 NAND2_X1 _19852_ (.A1(_07095_),
    .A2(_07795_),
    .ZN(_10192_));
 NAND2_X1 _19853_ (.A1(_07095_),
    .A2(_08365_),
    .ZN(_10193_));
 NAND4_X1 _19854_ (.A1(_10190_),
    .A2(_10191_),
    .A3(_10192_),
    .A4(_10193_),
    .ZN(_10194_));
 NAND2_X1 _19855_ (.A1(_08422_),
    .A2(_08167_),
    .ZN(_10195_));
 NAND4_X1 _19856_ (.A1(_08080_),
    .A2(_08478_),
    .A3(_07554_),
    .A4(_08403_),
    .ZN(_10196_));
 OAI211_X1 _19857_ (.A(_10195_),
    .B(_10196_),
    .C1(_07685_),
    .C2(_09310_),
    .ZN(_10197_));
 AOI21_X1 _19858_ (.A(_07685_),
    .B1(_09264_),
    .B2(_09484_),
    .ZN(_10198_));
 NOR2_X1 _19859_ (.A1(_07685_),
    .A2(_09347_),
    .ZN(_10199_));
 NOR4_X1 _19860_ (.A1(_10194_),
    .A2(_10197_),
    .A3(_10198_),
    .A4(_10199_),
    .ZN(_10200_));
 NAND2_X1 _19861_ (.A1(_08156_),
    .A2(_08308_),
    .ZN(_10201_));
 OAI211_X1 _19862_ (.A(_08178_),
    .B(_10201_),
    .C1(_09320_),
    .C2(_07707_),
    .ZN(_10202_));
 NAND4_X1 _19863_ (.A1(_08080_),
    .A2(_08478_),
    .A3(_07598_),
    .A4(_08113_),
    .ZN(_10203_));
 OAI211_X1 _19864_ (.A(_09309_),
    .B(_10203_),
    .C1(_07663_),
    .C2(_09311_),
    .ZN(_10204_));
 OAI21_X1 _19865_ (.A(_09869_),
    .B1(_09320_),
    .B2(_08482_),
    .ZN(_10205_));
 NOR4_X1 _19866_ (.A1(_10202_),
    .A2(_10204_),
    .A3(_10205_),
    .A4(_09317_),
    .ZN(_10206_));
 OAI21_X1 _19867_ (.A(_07839_),
    .B1(_07981_),
    .B2(_08233_),
    .ZN(_10207_));
 OAI211_X1 _19868_ (.A(_07411_),
    .B(_07194_),
    .C1(_08459_),
    .C2(_08102_),
    .ZN(_10208_));
 OAI21_X1 _19869_ (.A(_07411_),
    .B1(_07216_),
    .B2(_09456_),
    .ZN(_10209_));
 OAI211_X1 _19870_ (.A(_07839_),
    .B(_08431_),
    .C1(_08478_),
    .C2(_07194_),
    .ZN(_10210_));
 AND4_X1 _19871_ (.A1(_10207_),
    .A2(_10208_),
    .A3(_10209_),
    .A4(_10210_),
    .ZN(_10211_));
 NAND4_X1 _19872_ (.A1(_10189_),
    .A2(_10200_),
    .A3(_10206_),
    .A4(_10211_),
    .ZN(_10212_));
 AOI21_X1 _19873_ (.A(_09468_),
    .B1(_09349_),
    .B2(_09314_),
    .ZN(_10213_));
 NAND2_X1 _19874_ (.A1(_07631_),
    .A2(_09321_),
    .ZN(_10214_));
 OAI211_X1 _19875_ (.A(_09363_),
    .B(_10214_),
    .C1(_09364_),
    .C2(_08102_),
    .ZN(_10215_));
 NOR2_X1 _19876_ (.A1(_08494_),
    .A2(_09468_),
    .ZN(_10216_));
 NOR4_X1 _19877_ (.A1(_08489_),
    .A2(_10213_),
    .A3(_10215_),
    .A4(_10216_),
    .ZN(_10217_));
 AND2_X1 _19878_ (.A1(_09489_),
    .A2(_09490_),
    .ZN(_10218_));
 NAND3_X1 _19879_ (.A1(_07784_),
    .A2(_08189_),
    .A3(_07543_),
    .ZN(_10219_));
 NAND3_X1 _19880_ (.A1(_07762_),
    .A2(_08189_),
    .A3(_07543_),
    .ZN(_10220_));
 NAND2_X1 _19881_ (.A1(_10219_),
    .A2(_10220_),
    .ZN(_10221_));
 AND2_X1 _19882_ (.A1(_08491_),
    .A2(_07904_),
    .ZN(_10222_));
 NOR2_X1 _19883_ (.A1(_10221_),
    .A2(_10222_),
    .ZN(_10223_));
 AND2_X1 _19884_ (.A1(_07194_),
    .A2(_07161_),
    .ZN(_10224_));
 OAI21_X1 _19885_ (.A(_07249_),
    .B1(_10224_),
    .B2(_07904_),
    .ZN(_10225_));
 OAI21_X1 _19886_ (.A(_08491_),
    .B1(_07861_),
    .B2(_09456_),
    .ZN(_10226_));
 AND4_X1 _19887_ (.A1(_10218_),
    .A2(_10223_),
    .A3(_10225_),
    .A4(_10226_),
    .ZN(_10227_));
 OAI21_X1 _19888_ (.A(_08450_),
    .B1(_08498_),
    .B2(_08473_),
    .ZN(_10228_));
 OAI21_X1 _19889_ (.A(_08450_),
    .B1(_09330_),
    .B2(_08455_),
    .ZN(_10229_));
 OAI211_X1 _19890_ (.A(_07576_),
    .B(_16714_),
    .C1(_16713_),
    .C2(_06875_),
    .ZN(_10230_));
 AND4_X1 _19891_ (.A1(_08472_),
    .A2(_10228_),
    .A3(_10229_),
    .A4(_10230_),
    .ZN(_10231_));
 OAI21_X1 _19892_ (.A(_07466_),
    .B1(_08413_),
    .B2(_09289_),
    .ZN(_10232_));
 OAI21_X1 _19893_ (.A(_09352_),
    .B1(_07795_),
    .B2(_08451_),
    .ZN(_10233_));
 OAI21_X1 _19894_ (.A(_09352_),
    .B1(_09324_),
    .B2(_09289_),
    .ZN(_10234_));
 AND4_X1 _19895_ (.A1(_09344_),
    .A2(_10232_),
    .A3(_10233_),
    .A4(_10234_),
    .ZN(_10235_));
 NAND4_X1 _19896_ (.A1(_10217_),
    .A2(_10227_),
    .A3(_10231_),
    .A4(_10235_),
    .ZN(_10236_));
 NOR2_X2 _19897_ (.A1(_10212_),
    .A2(_10236_),
    .ZN(_10237_));
 XOR2_X2 _19898_ (.A(_10181_),
    .B(_10237_),
    .Z(_10238_));
 XNOR2_X1 _19899_ (.A(_10120_),
    .B(_10238_),
    .ZN(_10239_));
 NAND3_X1 _19900_ (.A1(_08830_),
    .A2(_09029_),
    .A3(_08858_),
    .ZN(_10240_));
 NAND2_X1 _19901_ (.A1(_08847_),
    .A2(_08998_),
    .ZN(_10241_));
 NAND3_X1 _19902_ (.A1(_09009_),
    .A2(_08833_),
    .A3(_08825_),
    .ZN(_10242_));
 OR2_X1 _19903_ (.A1(_09057_),
    .A2(_09098_),
    .ZN(_10243_));
 AND4_X1 _19904_ (.A1(_10241_),
    .A2(_09071_),
    .A3(_10242_),
    .A4(_10243_),
    .ZN(_10244_));
 OAI21_X1 _19905_ (.A(_08830_),
    .B1(_09074_),
    .B2(_08889_),
    .ZN(_10245_));
 OAI211_X1 _19906_ (.A(_08829_),
    .B(_08843_),
    .C1(_08964_),
    .C2(_09115_),
    .ZN(_10246_));
 AND4_X1 _19907_ (.A1(_10240_),
    .A2(_10244_),
    .A3(_10245_),
    .A4(_10246_),
    .ZN(_10247_));
 NAND2_X1 _19908_ (.A1(_09106_),
    .A2(_09093_),
    .ZN(_10248_));
 OAI211_X1 _19909_ (.A(_08913_),
    .B(_08914_),
    .C1(_08882_),
    .C2(_08909_),
    .ZN(_10249_));
 AND4_X1 _19910_ (.A1(_10248_),
    .A2(_10249_),
    .A3(_09693_),
    .A4(_09928_),
    .ZN(_10250_));
 AND2_X1 _19911_ (.A1(_08874_),
    .A2(_08844_),
    .ZN(_10251_));
 OAI21_X1 _19912_ (.A(_09720_),
    .B1(_08882_),
    .B2(_10251_),
    .ZN(_10252_));
 OAI21_X1 _19913_ (.A(_09720_),
    .B1(_09074_),
    .B2(_09710_),
    .ZN(_10253_));
 AND3_X1 _19914_ (.A1(_10250_),
    .A2(_10252_),
    .A3(_10253_),
    .ZN(_10254_));
 NAND3_X1 _19915_ (.A1(_08860_),
    .A2(_08833_),
    .A3(_08914_),
    .ZN(_10255_));
 OAI21_X1 _19916_ (.A(_10255_),
    .B1(_08932_),
    .B2(_09142_),
    .ZN(_10256_));
 AOI21_X1 _19917_ (.A(_10256_),
    .B1(_08855_),
    .B2(_08936_),
    .ZN(_10257_));
 OAI211_X1 _19918_ (.A(_08940_),
    .B(_08868_),
    .C1(_08844_),
    .C2(_08878_),
    .ZN(_10258_));
 OAI21_X1 _19919_ (.A(_08940_),
    .B1(_08907_),
    .B2(_08894_),
    .ZN(_10259_));
 AND3_X1 _19920_ (.A1(_10258_),
    .A2(_10259_),
    .A3(_09708_),
    .ZN(_10260_));
 OAI21_X1 _19921_ (.A(_08936_),
    .B1(_08904_),
    .B2(_08853_),
    .ZN(_10261_));
 OAI21_X1 _19922_ (.A(_08936_),
    .B1(_09077_),
    .B2(_09710_),
    .ZN(_10262_));
 AND4_X1 _19923_ (.A1(_10257_),
    .A2(_10260_),
    .A3(_10261_),
    .A4(_10262_),
    .ZN(_10263_));
 OAI21_X1 _19924_ (.A(_09075_),
    .B1(_08943_),
    .B2(_09077_),
    .ZN(_10264_));
 NAND3_X1 _19925_ (.A1(_08821_),
    .A2(_08888_),
    .A3(_08824_),
    .ZN(_10265_));
 NAND2_X1 _19926_ (.A1(_09009_),
    .A2(_08888_),
    .ZN(_10266_));
 AND4_X1 _19927_ (.A1(_08883_),
    .A2(_10264_),
    .A3(_10265_),
    .A4(_10266_),
    .ZN(_10267_));
 NAND4_X1 _19928_ (.A1(_10247_),
    .A2(_10254_),
    .A3(_10263_),
    .A4(_10267_),
    .ZN(_10268_));
 NAND4_X1 _19929_ (.A1(_09003_),
    .A2(_08973_),
    .A3(_08886_),
    .A4(_08868_),
    .ZN(_10269_));
 NAND2_X1 _19930_ (.A1(_09975_),
    .A2(_09051_),
    .ZN(_10270_));
 AND2_X1 _19931_ (.A1(_09026_),
    .A2(_08903_),
    .ZN(_10271_));
 AND2_X1 _19932_ (.A1(_09025_),
    .A2(_08859_),
    .ZN(_10272_));
 NOR4_X1 _19933_ (.A1(_10270_),
    .A2(_10271_),
    .A3(_10272_),
    .A4(_09699_),
    .ZN(_10273_));
 OAI211_X1 _19934_ (.A(_09031_),
    .B(_09107_),
    .C1(_08844_),
    .C2(_08878_),
    .ZN(_10274_));
 AND4_X1 _19935_ (.A1(_08878_),
    .A2(_09003_),
    .A3(_08886_),
    .A4(_08842_),
    .ZN(_10275_));
 AND2_X1 _19936_ (.A1(_09020_),
    .A2(_08855_),
    .ZN(_10276_));
 AOI221_X1 _19937_ (.A(_10275_),
    .B1(_09925_),
    .B2(_09020_),
    .C1(_08973_),
    .C2(_10276_),
    .ZN(_10277_));
 AND4_X1 _19938_ (.A1(_10269_),
    .A2(_10273_),
    .A3(_10274_),
    .A4(_10277_),
    .ZN(_10278_));
 OAI211_X1 _19939_ (.A(_08993_),
    .B(_09107_),
    .C1(_08964_),
    .C2(_08858_),
    .ZN(_10279_));
 OAI211_X1 _19940_ (.A(_08993_),
    .B(_08874_),
    .C1(_08973_),
    .C2(_08878_),
    .ZN(_10280_));
 OAI21_X1 _19941_ (.A(_08994_),
    .B1(_08965_),
    .B2(_08915_),
    .ZN(_10281_));
 AND4_X1 _19942_ (.A1(_09141_),
    .A2(_10279_),
    .A3(_10280_),
    .A4(_10281_),
    .ZN(_10282_));
 OAI21_X1 _19943_ (.A(_08957_),
    .B1(_09014_),
    .B2(_08836_),
    .ZN(_10283_));
 OAI21_X1 _19944_ (.A(_10283_),
    .B1(_09056_),
    .B2(_09143_),
    .ZN(_10284_));
 NAND2_X1 _19945_ (.A1(_08969_),
    .A2(_08957_),
    .ZN(_10285_));
 NAND2_X1 _19946_ (.A1(_08960_),
    .A2(_10285_),
    .ZN(_10286_));
 NOR4_X1 _19947_ (.A1(_10284_),
    .A2(_10286_),
    .A3(_09124_),
    .A4(_08961_),
    .ZN(_10287_));
 OAI21_X1 _19948_ (.A(_08982_),
    .B1(_08943_),
    .B2(_08838_),
    .ZN(_10288_));
 OAI21_X1 _19949_ (.A(_08976_),
    .B1(_08933_),
    .B2(_08923_),
    .ZN(_10289_));
 OAI21_X1 _19950_ (.A(_08976_),
    .B1(_08969_),
    .B2(_08850_),
    .ZN(_10290_));
 OAI211_X1 _19951_ (.A(_08913_),
    .B(_08950_),
    .C1(_08908_),
    .C2(_09009_),
    .ZN(_10291_));
 AND4_X1 _19952_ (.A1(_10288_),
    .A2(_10289_),
    .A3(_10290_),
    .A4(_10291_),
    .ZN(_10292_));
 NAND3_X1 _19953_ (.A1(_08821_),
    .A2(_08824_),
    .A3(_08951_),
    .ZN(_10293_));
 NAND2_X1 _19954_ (.A1(_08952_),
    .A2(_08909_),
    .ZN(_10294_));
 NAND2_X1 _19955_ (.A1(_08943_),
    .A2(_08952_),
    .ZN(_10295_));
 AND4_X1 _19956_ (.A1(_08971_),
    .A2(_10293_),
    .A3(_10294_),
    .A4(_10295_),
    .ZN(_10296_));
 AND4_X1 _19957_ (.A1(_10282_),
    .A2(_10287_),
    .A3(_10292_),
    .A4(_10296_),
    .ZN(_10297_));
 NOR2_X1 _19958_ (.A1(_09109_),
    .A2(_09916_),
    .ZN(_10298_));
 INV_X1 _19959_ (.A(_09095_),
    .ZN(_10299_));
 AOI21_X1 _19960_ (.A(_09109_),
    .B1(_10299_),
    .B2(_08893_),
    .ZN(_10300_));
 AOI211_X1 _19961_ (.A(_10298_),
    .B(_10300_),
    .C1(_09050_),
    .C2(_09005_),
    .ZN(_10301_));
 AND2_X1 _19962_ (.A1(_08938_),
    .A2(_09008_),
    .ZN(_10302_));
 AND2_X1 _19963_ (.A1(_09007_),
    .A2(_08843_),
    .ZN(_10303_));
 AND2_X1 _19964_ (.A1(_09007_),
    .A2(_09077_),
    .ZN(_10304_));
 NOR4_X1 _19965_ (.A1(_10302_),
    .A2(_10303_),
    .A3(_09959_),
    .A4(_10304_),
    .ZN(_10305_));
 NAND4_X1 _19966_ (.A1(_10278_),
    .A2(_10297_),
    .A3(_10301_),
    .A4(_10305_),
    .ZN(_10306_));
 NOR2_X2 _19967_ (.A1(_10268_),
    .A2(_10306_),
    .ZN(_10307_));
 XOR2_X2 _19968_ (.A(_10307_),
    .B(_09035_),
    .Z(_10308_));
 XNOR2_X1 _19969_ (.A(_10239_),
    .B(_10308_),
    .ZN(_10309_));
 XNOR2_X1 _19970_ (.A(_10309_),
    .B(_17093_),
    .ZN(_10310_));
 MUX2_X1 _19971_ (.A(_10064_),
    .B(_10310_),
    .S(_09040_),
    .Z(_00728_));
 XOR2_X1 _19972_ (.A(_17094_),
    .B(_17018_),
    .Z(_10311_));
 AND2_X1 _19973_ (.A1(_04340_),
    .A2(_05390_),
    .ZN(_10312_));
 OR2_X1 _19974_ (.A1(_05467_),
    .A2(_10312_),
    .ZN(_10313_));
 NAND2_X1 _19975_ (.A1(_06116_),
    .A2(_05401_),
    .ZN(_10314_));
 OAI21_X1 _19976_ (.A(_10314_),
    .B1(_05423_),
    .B2(_09183_),
    .ZN(_10315_));
 AOI21_X1 _19977_ (.A(_05423_),
    .B1(_09200_),
    .B2(_09185_),
    .ZN(_10316_));
 OR4_X1 _19978_ (.A1(_09151_),
    .A2(_10313_),
    .A3(_10315_),
    .A4(_10316_),
    .ZN(_10317_));
 OAI211_X1 _19979_ (.A(_05522_),
    .B(_05863_),
    .C1(_06314_),
    .C2(_06325_),
    .ZN(_10318_));
 OAI21_X1 _19980_ (.A(_05522_),
    .B1(_05096_),
    .B2(_06490_),
    .ZN(_10319_));
 OAI211_X1 _19981_ (.A(_10318_),
    .B(_10319_),
    .C1(_05918_),
    .C2(_09168_),
    .ZN(_10320_));
 AND3_X1 _19982_ (.A1(_05445_),
    .A2(_05687_),
    .A3(_05324_),
    .ZN(_10321_));
 OR3_X1 _19983_ (.A1(_10056_),
    .A2(_09162_),
    .A3(_10321_),
    .ZN(_10322_));
 AND2_X1 _19984_ (.A1(_05258_),
    .A2(_05445_),
    .ZN(_10323_));
 INV_X1 _19985_ (.A(_10323_),
    .ZN(_10324_));
 AND4_X1 _19986_ (.A1(_09176_),
    .A2(_10324_),
    .A3(_09641_),
    .A4(_10099_),
    .ZN(_10325_));
 INV_X1 _19987_ (.A(_09173_),
    .ZN(_10326_));
 AND2_X1 _19988_ (.A1(_05291_),
    .A2(_05159_),
    .ZN(_10327_));
 INV_X1 _19989_ (.A(_10327_),
    .ZN(_10328_));
 NAND4_X1 _19990_ (.A1(_10325_),
    .A2(_10326_),
    .A3(_10029_),
    .A4(_10328_),
    .ZN(_10329_));
 NOR4_X1 _19991_ (.A1(_10317_),
    .A2(_10320_),
    .A3(_10322_),
    .A4(_10329_),
    .ZN(_10330_));
 NOR4_X1 _19992_ (.A1(_10078_),
    .A2(_09211_),
    .A3(_09212_),
    .A4(_09213_),
    .ZN(_10331_));
 AND2_X1 _19993_ (.A1(_05676_),
    .A2(_06556_),
    .ZN(_10332_));
 AND2_X1 _19994_ (.A1(_04559_),
    .A2(_06556_),
    .ZN(_10333_));
 AND2_X1 _19995_ (.A1(_04625_),
    .A2(_06545_),
    .ZN(_10334_));
 NOR4_X1 _19996_ (.A1(_10332_),
    .A2(_10333_),
    .A3(_10066_),
    .A4(_10334_),
    .ZN(_10335_));
 OAI21_X1 _19997_ (.A(_06391_),
    .B1(_10008_),
    .B2(_04669_),
    .ZN(_10336_));
 AND4_X1 _19998_ (.A1(_09221_),
    .A2(_10335_),
    .A3(_09681_),
    .A4(_10336_),
    .ZN(_10337_));
 OAI221_X1 _19999_ (.A(_06281_),
    .B1(_06314_),
    .B2(_05203_),
    .C1(_05863_),
    .C2(_05797_),
    .ZN(_10338_));
 AOI21_X1 _20000_ (.A(_06215_),
    .B1(_06127_),
    .B2(_09183_),
    .ZN(_10339_));
 OAI22_X1 _20001_ (.A1(_10075_),
    .A2(_05313_),
    .B1(_06215_),
    .B2(_05918_),
    .ZN(_10340_));
 AOI211_X1 _20002_ (.A(_10339_),
    .B(_10340_),
    .C1(_06171_),
    .C2(_09639_),
    .ZN(_10341_));
 AND4_X1 _20003_ (.A1(_10331_),
    .A2(_10337_),
    .A3(_10338_),
    .A4(_10341_),
    .ZN(_10342_));
 NAND4_X1 _20004_ (.A1(_04461_),
    .A2(_09158_),
    .A3(_04959_),
    .A4(_06303_),
    .ZN(_10343_));
 NAND3_X1 _20005_ (.A1(_04263_),
    .A2(_04461_),
    .A3(_05687_),
    .ZN(_10344_));
 AND3_X1 _20006_ (.A1(_05036_),
    .A2(_10343_),
    .A3(_10344_),
    .ZN(_10345_));
 OAI21_X1 _20007_ (.A(_05045_),
    .B1(_06116_),
    .B2(_09182_),
    .ZN(_10346_));
 OAI21_X1 _20008_ (.A(_04614_),
    .B1(_05676_),
    .B2(_04855_),
    .ZN(_10347_));
 NAND4_X1 _20009_ (.A1(_10345_),
    .A2(_04702_),
    .A3(_10346_),
    .A4(_10347_),
    .ZN(_10348_));
 NAND2_X1 _20010_ (.A1(_04209_),
    .A2(_05225_),
    .ZN(_10349_));
 OAI21_X1 _20011_ (.A(_04494_),
    .B1(_05082_),
    .B2(_05962_),
    .ZN(_10350_));
 NAND4_X1 _20012_ (.A1(_04285_),
    .A2(_10349_),
    .A3(_09666_),
    .A4(_10350_),
    .ZN(_10351_));
 OAI21_X1 _20013_ (.A(_10087_),
    .B1(_09193_),
    .B2(_05126_),
    .ZN(_10352_));
 NAND3_X1 _20014_ (.A1(_04931_),
    .A2(_04940_),
    .A3(_09661_),
    .ZN(_10353_));
 NOR4_X1 _20015_ (.A1(_10348_),
    .A2(_10351_),
    .A3(_10352_),
    .A4(_10353_),
    .ZN(_10354_));
 AND2_X1 _20016_ (.A1(_04340_),
    .A2(_06017_),
    .ZN(_10355_));
 INV_X1 _20017_ (.A(_10355_),
    .ZN(_10356_));
 AND3_X1 _20018_ (.A1(_09245_),
    .A2(_10356_),
    .A3(_06061_),
    .ZN(_10357_));
 OAI21_X1 _20019_ (.A(_09251_),
    .B1(_04559_),
    .B2(_04395_),
    .ZN(_10358_));
 OAI21_X1 _20020_ (.A(_09251_),
    .B1(_04746_),
    .B2(_04778_),
    .ZN(_10359_));
 OAI21_X1 _20021_ (.A(_09246_),
    .B1(_05599_),
    .B2(_10008_),
    .ZN(_10360_));
 NAND4_X1 _20022_ (.A1(_10357_),
    .A2(_10358_),
    .A3(_10359_),
    .A4(_10360_),
    .ZN(_10361_));
 OAI21_X1 _20023_ (.A(_05786_),
    .B1(_09623_),
    .B2(_10011_),
    .ZN(_10362_));
 NAND4_X1 _20024_ (.A1(_05786_),
    .A2(_06303_),
    .A3(_04899_),
    .A4(_06236_),
    .ZN(_10363_));
 OAI211_X1 _20025_ (.A(_10362_),
    .B(_10363_),
    .C1(_06402_),
    .C2(_09238_),
    .ZN(_10364_));
 AND2_X1 _20026_ (.A1(_05632_),
    .A2(_04263_),
    .ZN(_10365_));
 INV_X1 _20027_ (.A(_10365_),
    .ZN(_10366_));
 OAI211_X1 _20028_ (.A(_10366_),
    .B(_09621_),
    .C1(_05434_),
    .C2(_05654_),
    .ZN(_10367_));
 OAI21_X1 _20029_ (.A(_05643_),
    .B1(_05654_),
    .B2(_04526_),
    .ZN(_10368_));
 NOR4_X1 _20030_ (.A1(_10361_),
    .A2(_10364_),
    .A3(_10367_),
    .A4(_10368_),
    .ZN(_10369_));
 NAND4_X1 _20031_ (.A1(_10330_),
    .A2(_10342_),
    .A3(_10354_),
    .A4(_10369_),
    .ZN(_10370_));
 NOR2_X2 _20032_ (.A1(_10370_),
    .A2(_06672_),
    .ZN(_10371_));
 XNOR2_X1 _20033_ (.A(_10371_),
    .B(_10181_),
    .ZN(_10372_));
 INV_X1 _20034_ (.A(_07400_),
    .ZN(_10373_));
 AOI21_X1 _20035_ (.A(_10373_),
    .B1(_09264_),
    .B2(_09484_),
    .ZN(_10374_));
 AND2_X1 _20036_ (.A1(_07948_),
    .A2(_07400_),
    .ZN(_10375_));
 AND4_X1 _20037_ (.A1(_08478_),
    .A2(_07150_),
    .A3(_07554_),
    .A4(_08463_),
    .ZN(_10376_));
 NOR3_X1 _20038_ (.A1(_10374_),
    .A2(_10375_),
    .A3(_10376_),
    .ZN(_10377_));
 AND2_X1 _20039_ (.A1(_08025_),
    .A2(_08451_),
    .ZN(_10378_));
 AOI21_X1 _20040_ (.A(_09292_),
    .B1(_08468_),
    .B2(_07282_),
    .ZN(_10379_));
 AOI211_X1 _20041_ (.A(_10378_),
    .B(_10379_),
    .C1(_08025_),
    .C2(_09887_),
    .ZN(_10380_));
 OAI221_X1 _20042_ (.A(_06732_),
    .B1(_06754_),
    .B2(_07161_),
    .C1(_08069_),
    .C2(_08233_),
    .ZN(_10381_));
 AND3_X1 _20043_ (.A1(_10381_),
    .A2(_09525_),
    .A3(_09297_),
    .ZN(_10382_));
 INV_X1 _20044_ (.A(_09530_),
    .ZN(_10383_));
 AND2_X1 _20045_ (.A1(_07356_),
    .A2(_06853_),
    .ZN(_10384_));
 INV_X1 _20046_ (.A(_10384_),
    .ZN(_10385_));
 AOI21_X1 _20047_ (.A(_09304_),
    .B1(_10385_),
    .B2(_07128_),
    .ZN(_10386_));
 AOI211_X1 _20048_ (.A(_10383_),
    .B(_10386_),
    .C1(_07839_),
    .C2(_09296_),
    .ZN(_10387_));
 AND4_X1 _20049_ (.A1(_10377_),
    .A2(_10380_),
    .A3(_10382_),
    .A4(_10387_),
    .ZN(_10388_));
 AND3_X1 _20050_ (.A1(_07784_),
    .A2(_08189_),
    .A3(_07062_),
    .ZN(_10389_));
 AOI211_X1 _20051_ (.A(_10389_),
    .B(_09499_),
    .C1(_06952_),
    .C2(_08156_),
    .ZN(_10390_));
 NAND4_X1 _20052_ (.A1(_08200_),
    .A2(_08461_),
    .A3(_08080_),
    .A4(_08403_),
    .ZN(_10391_));
 AND3_X1 _20053_ (.A1(_10390_),
    .A2(_09869_),
    .A3(_10391_),
    .ZN(_10392_));
 OAI21_X1 _20054_ (.A(_07893_),
    .B1(_07762_),
    .B2(_08498_),
    .ZN(_10393_));
 AND3_X1 _20055_ (.A1(_10393_),
    .A2(_08124_),
    .A3(_08058_),
    .ZN(_10394_));
 AND2_X1 _20056_ (.A1(_07084_),
    .A2(_07795_),
    .ZN(_10395_));
 AOI211_X1 _20057_ (.A(_09843_),
    .B(_10395_),
    .C1(_07095_),
    .C2(_08473_),
    .ZN(_10396_));
 OAI21_X1 _20058_ (.A(_08422_),
    .B1(_07532_),
    .B2(_08167_),
    .ZN(_10397_));
 AND4_X1 _20059_ (.A1(_08441_),
    .A2(_09514_),
    .A3(_08447_),
    .A4(_10397_),
    .ZN(_10398_));
 AND4_X1 _20060_ (.A1(_10392_),
    .A2(_10394_),
    .A3(_10396_),
    .A4(_10398_),
    .ZN(_10399_));
 AND4_X1 _20061_ (.A1(_07150_),
    .A2(_08211_),
    .A3(_07183_),
    .A4(_06974_),
    .ZN(_10400_));
 AND2_X1 _20062_ (.A1(_07631_),
    .A2(_07762_),
    .ZN(_10401_));
 AOI211_X1 _20063_ (.A(_10400_),
    .B(_10401_),
    .C1(_08485_),
    .C2(_07904_),
    .ZN(_10402_));
 INV_X1 _20064_ (.A(_07337_),
    .ZN(_10403_));
 NAND2_X1 _20065_ (.A1(_09277_),
    .A2(_10403_),
    .ZN(_10404_));
 OAI21_X1 _20066_ (.A(_07466_),
    .B1(_10404_),
    .B2(_07861_),
    .ZN(_10405_));
 OAI211_X1 _20067_ (.A(_08189_),
    .B(_08222_),
    .C1(_06952_),
    .C2(_07029_),
    .ZN(_10406_));
 AND4_X1 _20068_ (.A1(_09461_),
    .A2(_09878_),
    .A3(_10405_),
    .A4(_10406_),
    .ZN(_10407_));
 OAI211_X1 _20069_ (.A(_06974_),
    .B(_08222_),
    .C1(_09289_),
    .C2(_09456_),
    .ZN(_10408_));
 AOI21_X1 _20070_ (.A(_09468_),
    .B1(_09287_),
    .B2(_07970_),
    .ZN(_10409_));
 NAND2_X1 _20071_ (.A1(_07315_),
    .A2(_07378_),
    .ZN(_10410_));
 OAI21_X1 _20072_ (.A(_10410_),
    .B1(_09468_),
    .B2(_08482_),
    .ZN(_10411_));
 AND2_X1 _20073_ (.A1(_07315_),
    .A2(_09321_),
    .ZN(_10412_));
 NOR4_X1 _20074_ (.A1(_10409_),
    .A2(_10411_),
    .A3(_06897_),
    .A4(_10412_),
    .ZN(_10413_));
 AND4_X1 _20075_ (.A1(_10402_),
    .A2(_10407_),
    .A3(_10408_),
    .A4(_10413_),
    .ZN(_10414_));
 AND2_X1 _20076_ (.A1(_07238_),
    .A2(_07904_),
    .ZN(_10415_));
 AND4_X1 _20077_ (.A1(_07194_),
    .A2(_07238_),
    .A3(_07850_),
    .A4(_08431_),
    .ZN(_10416_));
 AOI211_X1 _20078_ (.A(_10415_),
    .B(_10416_),
    .C1(_07249_),
    .C2(_06776_),
    .ZN(_10417_));
 OAI21_X1 _20079_ (.A(_08450_),
    .B1(_07652_),
    .B2(_07904_),
    .ZN(_10418_));
 AND3_X1 _20080_ (.A1(_07565_),
    .A2(_07183_),
    .A3(_07598_),
    .ZN(_10419_));
 AOI211_X1 _20081_ (.A(_10419_),
    .B(_09260_),
    .C1(_07532_),
    .C2(_07576_),
    .ZN(_10420_));
 OAI21_X1 _20082_ (.A(_07007_),
    .B1(_08047_),
    .B2(_07948_),
    .ZN(_10421_));
 OAI21_X1 _20083_ (.A(_07576_),
    .B1(_09327_),
    .B2(_10384_),
    .ZN(_10422_));
 AND4_X1 _20084_ (.A1(_10418_),
    .A2(_10420_),
    .A3(_10421_),
    .A4(_10422_),
    .ZN(_10423_));
 OAI21_X1 _20085_ (.A(_07249_),
    .B1(_09313_),
    .B2(_09837_),
    .ZN(_10424_));
 NAND3_X1 _20086_ (.A1(_06776_),
    .A2(_08200_),
    .A3(_07543_),
    .ZN(_10425_));
 INV_X1 _20087_ (.A(_10222_),
    .ZN(_10426_));
 OAI21_X1 _20088_ (.A(_08491_),
    .B1(_09330_),
    .B2(_07948_),
    .ZN(_10427_));
 AND4_X1 _20089_ (.A1(_10425_),
    .A2(_10426_),
    .A3(_10219_),
    .A4(_10427_),
    .ZN(_10428_));
 AND4_X1 _20090_ (.A1(_10417_),
    .A2(_10423_),
    .A3(_10424_),
    .A4(_10428_),
    .ZN(_10429_));
 NAND4_X1 _20091_ (.A1(_10388_),
    .A2(_10399_),
    .A3(_10414_),
    .A4(_10429_),
    .ZN(_10430_));
 NOR2_X2 _20092_ (.A1(_10430_),
    .A2(_07040_),
    .ZN(_10431_));
 OAI21_X1 _20093_ (.A(_08592_),
    .B1(_08698_),
    .B2(_09810_),
    .ZN(_10432_));
 OAI21_X1 _20094_ (.A(_08592_),
    .B1(_08601_),
    .B2(_08724_),
    .ZN(_10433_));
 NAND4_X1 _20095_ (.A1(_08592_),
    .A2(_08590_),
    .A3(_08587_),
    .A4(_08615_),
    .ZN(_10434_));
 AND3_X1 _20096_ (.A1(_10432_),
    .A2(_10433_),
    .A3(_10434_),
    .ZN(_10435_));
 OAI21_X1 _20097_ (.A(_08676_),
    .B1(_08519_),
    .B2(_08724_),
    .ZN(_10436_));
 AND3_X1 _20098_ (.A1(_08522_),
    .A2(_08509_),
    .A3(_08517_),
    .ZN(_10437_));
 AND2_X1 _20099_ (.A1(_08688_),
    .A2(_08523_),
    .ZN(_10438_));
 AOI211_X1 _20100_ (.A(_10437_),
    .B(_10438_),
    .C1(_08685_),
    .C2(_08523_),
    .ZN(_10439_));
 OAI21_X1 _20101_ (.A(_08676_),
    .B1(_08510_),
    .B2(_08568_),
    .ZN(_10440_));
 OAI21_X1 _20102_ (.A(_08523_),
    .B1(_08764_),
    .B2(_08661_),
    .ZN(_10441_));
 AND4_X1 _20103_ (.A1(_10436_),
    .A2(_10439_),
    .A3(_10440_),
    .A4(_10441_),
    .ZN(_10442_));
 AND2_X1 _20104_ (.A1(_08702_),
    .A2(_08724_),
    .ZN(_10443_));
 AND2_X1 _20105_ (.A1(_08714_),
    .A2(_08702_),
    .ZN(_10444_));
 AOI211_X1 _20106_ (.A(_10443_),
    .B(_10444_),
    .C1(_08703_),
    .C2(_08601_),
    .ZN(_10445_));
 OAI211_X1 _20107_ (.A(_08703_),
    .B(_08733_),
    .C1(_09382_),
    .C2(_08574_),
    .ZN(_10446_));
 AND4_X1 _20108_ (.A1(_10435_),
    .A2(_10442_),
    .A3(_10445_),
    .A4(_10446_),
    .ZN(_10447_));
 AND2_X1 _20109_ (.A1(_08663_),
    .A2(_08552_),
    .ZN(_10448_));
 AOI211_X1 _20110_ (.A(_10448_),
    .B(_08782_),
    .C1(_08663_),
    .C2(_08684_),
    .ZN(_10449_));
 OAI211_X1 _20111_ (.A(_08663_),
    .B(_08733_),
    .C1(_08651_),
    .C2(_08794_),
    .ZN(_10450_));
 OAI21_X1 _20112_ (.A(_08629_),
    .B1(_08594_),
    .B2(_08544_),
    .ZN(_10451_));
 AND4_X1 _20113_ (.A1(_08635_),
    .A2(_10449_),
    .A3(_10450_),
    .A4(_10451_),
    .ZN(_10452_));
 NAND3_X1 _20114_ (.A1(_08682_),
    .A2(_08632_),
    .A3(_08581_),
    .ZN(_10453_));
 AND4_X1 _20115_ (.A1(_09806_),
    .A2(_10122_),
    .A3(_10453_),
    .A4(_09808_),
    .ZN(_10454_));
 OAI21_X1 _20116_ (.A(_08549_),
    .B1(_08689_),
    .B2(_08621_),
    .ZN(_10455_));
 AND2_X1 _20117_ (.A1(_08510_),
    .A2(_08548_),
    .ZN(_10456_));
 AOI211_X1 _20118_ (.A(_10456_),
    .B(_08763_),
    .C1(_09548_),
    .C2(_08549_),
    .ZN(_10457_));
 AND4_X1 _20119_ (.A1(_10452_),
    .A2(_10454_),
    .A3(_10455_),
    .A4(_10457_),
    .ZN(_10458_));
 OAI21_X1 _20120_ (.A(_08541_),
    .B1(_09548_),
    .B2(_08531_),
    .ZN(_10459_));
 AOI21_X1 _20121_ (.A(_08788_),
    .B1(_08553_),
    .B2(_08541_),
    .ZN(_10460_));
 AND3_X1 _20122_ (.A1(_10141_),
    .A2(_09396_),
    .A3(_09397_),
    .ZN(_10461_));
 OAI221_X1 _20123_ (.A(_08622_),
    .B1(_08651_),
    .B2(_08507_),
    .C1(_08733_),
    .C2(_08637_),
    .ZN(_10462_));
 AND4_X1 _20124_ (.A1(_10459_),
    .A2(_10460_),
    .A3(_10461_),
    .A4(_10462_),
    .ZN(_10463_));
 OAI21_X1 _20125_ (.A(_08586_),
    .B1(_09404_),
    .B2(_08665_),
    .ZN(_10464_));
 AND2_X1 _20126_ (.A1(_08585_),
    .A2(_08707_),
    .ZN(_10465_));
 AOI211_X1 _20127_ (.A(_10465_),
    .B(_09541_),
    .C1(_08586_),
    .C2(_08661_),
    .ZN(_10466_));
 AND2_X1 _20128_ (.A1(_08510_),
    .A2(_08625_),
    .ZN(_10467_));
 AOI211_X1 _20129_ (.A(_08626_),
    .B(_10467_),
    .C1(_08637_),
    .C2(_08636_),
    .ZN(_10468_));
 AND4_X1 _20130_ (.A1(_10463_),
    .A2(_10464_),
    .A3(_10466_),
    .A4(_10468_),
    .ZN(_10469_));
 AND4_X1 _20131_ (.A1(_08618_),
    .A2(_08580_),
    .A3(_08563_),
    .A4(_08517_),
    .ZN(_10470_));
 AOI221_X4 _20132_ (.A(_10470_),
    .B1(_08724_),
    .B2(_08572_),
    .C1(_09436_),
    .C2(_08651_),
    .ZN(_10471_));
 INV_X1 _20133_ (.A(_09769_),
    .ZN(_10472_));
 NAND3_X1 _20134_ (.A1(_08553_),
    .A2(_08633_),
    .A3(_08641_),
    .ZN(_10473_));
 OAI21_X1 _20135_ (.A(_08650_),
    .B1(_08747_),
    .B2(_08667_),
    .ZN(_10474_));
 OAI21_X1 _20136_ (.A(_08604_),
    .B1(_08684_),
    .B2(_08679_),
    .ZN(_10475_));
 AND4_X1 _20137_ (.A1(_10472_),
    .A2(_10473_),
    .A3(_10474_),
    .A4(_10475_),
    .ZN(_10476_));
 OAI211_X1 _20138_ (.A(_08641_),
    .B(_08581_),
    .C1(_08708_),
    .C2(_08607_),
    .ZN(_10477_));
 NAND3_X1 _20139_ (.A1(_08708_),
    .A2(_08641_),
    .A3(_08642_),
    .ZN(_10478_));
 OAI21_X1 _20140_ (.A(_08609_),
    .B1(_08758_),
    .B2(_08611_),
    .ZN(_10479_));
 OAI21_X1 _20141_ (.A(_08609_),
    .B1(_08568_),
    .B2(_08797_),
    .ZN(_10480_));
 NAND3_X1 _20142_ (.A1(_08715_),
    .A2(_08641_),
    .A3(_08642_),
    .ZN(_10481_));
 AND4_X1 _20143_ (.A1(_10478_),
    .A2(_10479_),
    .A3(_10480_),
    .A4(_10481_),
    .ZN(_10482_));
 AND4_X1 _20144_ (.A1(_10471_),
    .A2(_10476_),
    .A3(_10477_),
    .A4(_10482_),
    .ZN(_10483_));
 NAND4_X1 _20145_ (.A1(_10447_),
    .A2(_10458_),
    .A3(_10469_),
    .A4(_10483_),
    .ZN(_10484_));
 NOR2_X2 _20146_ (.A1(_10484_),
    .A2(_08696_),
    .ZN(_10485_));
 XNOR2_X2 _20147_ (.A(_10431_),
    .B(_10485_),
    .ZN(_10486_));
 XNOR2_X1 _20148_ (.A(_10372_),
    .B(_10486_),
    .ZN(_10487_));
 AOI221_X4 _20149_ (.A(_09705_),
    .B1(_08911_),
    .B2(_09026_),
    .C1(_08844_),
    .C2(_09699_),
    .ZN(_10488_));
 OAI21_X1 _20150_ (.A(_09031_),
    .B1(_08986_),
    .B2(_08838_),
    .ZN(_10489_));
 OAI21_X1 _20151_ (.A(_09031_),
    .B1(_08938_),
    .B2(_08882_),
    .ZN(_10490_));
 AND4_X1 _20152_ (.A1(_09092_),
    .A2(_10488_),
    .A3(_10489_),
    .A4(_10490_),
    .ZN(_10491_));
 INV_X1 _20153_ (.A(_09077_),
    .ZN(_10492_));
 AOI21_X1 _20154_ (.A(_08983_),
    .B1(_10492_),
    .B2(_09111_),
    .ZN(_10493_));
 NAND3_X1 _20155_ (.A1(_09087_),
    .A2(_09029_),
    .A3(_08823_),
    .ZN(_10494_));
 NAND2_X1 _20156_ (.A1(_09087_),
    .A2(_08843_),
    .ZN(_10495_));
 OAI211_X1 _20157_ (.A(_10494_),
    .B(_10495_),
    .C1(_09056_),
    .C2(_08995_),
    .ZN(_10496_));
 NOR4_X1 _20158_ (.A1(_10493_),
    .A2(_10496_),
    .A3(_09951_),
    .A4(_09700_),
    .ZN(_10497_));
 OAI211_X1 _20159_ (.A(_08972_),
    .B(_09029_),
    .C1(_08973_),
    .C2(_08878_),
    .ZN(_10498_));
 OAI21_X1 _20160_ (.A(_08972_),
    .B1(_08838_),
    .B2(_08989_),
    .ZN(_10499_));
 NAND4_X1 _20161_ (.A1(_10498_),
    .A2(_10499_),
    .A3(_08955_),
    .A4(_10294_),
    .ZN(_10500_));
 AND2_X1 _20162_ (.A1(_09053_),
    .A2(_08836_),
    .ZN(_10501_));
 AND2_X1 _20163_ (.A1(_09690_),
    .A2(_09053_),
    .ZN(_10502_));
 NOR4_X1 _20164_ (.A1(_09966_),
    .A2(_10500_),
    .A3(_10501_),
    .A4(_10502_),
    .ZN(_10503_));
 AOI22_X1 _20165_ (.A1(_10303_),
    .A2(_09116_),
    .B1(_08853_),
    .B2(_09008_),
    .ZN(_10504_));
 OAI21_X1 _20166_ (.A(_09005_),
    .B1(_08919_),
    .B2(_08853_),
    .ZN(_10505_));
 OAI21_X1 _20167_ (.A(_09008_),
    .B1(_08954_),
    .B2(_09710_),
    .ZN(_10506_));
 AND4_X1 _20168_ (.A1(_09714_),
    .A2(_10504_),
    .A3(_10505_),
    .A4(_10506_),
    .ZN(_10507_));
 NAND4_X1 _20169_ (.A1(_10491_),
    .A2(_10497_),
    .A3(_10503_),
    .A4(_10507_),
    .ZN(_10508_));
 AND2_X1 _20170_ (.A1(_08901_),
    .A2(_08923_),
    .ZN(_10509_));
 AND2_X1 _20171_ (.A1(_08901_),
    .A2(_08965_),
    .ZN(_10510_));
 AOI211_X1 _20172_ (.A(_10509_),
    .B(_10510_),
    .C1(_08987_),
    .C2(_09720_),
    .ZN(_10511_));
 NAND2_X1 _20173_ (.A1(_09720_),
    .A2(_08843_),
    .ZN(_10512_));
 NAND2_X1 _20174_ (.A1(_09017_),
    .A2(_08906_),
    .ZN(_10513_));
 NAND2_X1 _20175_ (.A1(_08906_),
    .A2(_08954_),
    .ZN(_10514_));
 OAI211_X1 _20176_ (.A(_08906_),
    .B(_08843_),
    .C1(_08844_),
    .C2(_08845_),
    .ZN(_10515_));
 AND4_X1 _20177_ (.A1(_10248_),
    .A2(_10513_),
    .A3(_10514_),
    .A4(_10515_),
    .ZN(_10516_));
 AND4_X1 _20178_ (.A1(_08905_),
    .A2(_10511_),
    .A3(_10512_),
    .A4(_10516_),
    .ZN(_10517_));
 NAND2_X1 _20179_ (.A1(_08936_),
    .A2(_08989_),
    .ZN(_10518_));
 NAND2_X1 _20180_ (.A1(_08936_),
    .A2(_08987_),
    .ZN(_10519_));
 NAND3_X1 _20181_ (.A1(_08931_),
    .A2(_10518_),
    .A3(_10519_),
    .ZN(_10520_));
 AOI21_X1 _20182_ (.A(_08932_),
    .B1(_08893_),
    .B2(_09142_),
    .ZN(_10521_));
 NAND3_X1 _20183_ (.A1(_08954_),
    .A2(_08827_),
    .A3(_08914_),
    .ZN(_10522_));
 NAND3_X1 _20184_ (.A1(_09710_),
    .A2(_08827_),
    .A3(_08914_),
    .ZN(_10523_));
 NAND3_X1 _20185_ (.A1(_09136_),
    .A2(_10522_),
    .A3(_10523_),
    .ZN(_10524_));
 NOR4_X1 _20186_ (.A1(_10520_),
    .A2(_10521_),
    .A3(_10524_),
    .A4(_09733_),
    .ZN(_10525_));
 NAND3_X1 _20187_ (.A1(_08830_),
    .A2(_08964_),
    .A3(_09107_),
    .ZN(_10526_));
 NAND3_X1 _20188_ (.A1(_08830_),
    .A2(_09029_),
    .A3(_08964_),
    .ZN(_10527_));
 NAND2_X1 _20189_ (.A1(_09122_),
    .A2(_08830_),
    .ZN(_10528_));
 NAND4_X1 _20190_ (.A1(_09942_),
    .A2(_10526_),
    .A3(_10527_),
    .A4(_10528_),
    .ZN(_10529_));
 AND2_X1 _20191_ (.A1(_08847_),
    .A2(_09710_),
    .ZN(_10530_));
 AOI21_X1 _20192_ (.A(_09057_),
    .B1(_08996_),
    .B2(_08895_),
    .ZN(_10531_));
 NOR4_X1 _20193_ (.A1(_10529_),
    .A2(_08839_),
    .A3(_10530_),
    .A4(_10531_),
    .ZN(_10532_));
 INV_X1 _20194_ (.A(_09073_),
    .ZN(_10533_));
 NAND2_X1 _20195_ (.A1(_09075_),
    .A2(_08855_),
    .ZN(_10534_));
 NAND3_X1 _20196_ (.A1(_09075_),
    .A2(_08824_),
    .A3(_09118_),
    .ZN(_10535_));
 NAND3_X1 _20197_ (.A1(_10533_),
    .A2(_10534_),
    .A3(_10535_),
    .ZN(_10536_));
 OAI21_X1 _20198_ (.A(_08888_),
    .B1(_08907_),
    .B2(_08909_),
    .ZN(_10537_));
 NAND4_X1 _20199_ (.A1(_09107_),
    .A2(_08886_),
    .A3(_08858_),
    .A4(_08825_),
    .ZN(_10538_));
 OAI211_X1 _20200_ (.A(_10537_),
    .B(_10538_),
    .C1(_08892_),
    .C2(_08999_),
    .ZN(_10539_));
 NOR4_X1 _20201_ (.A1(_10536_),
    .A2(_10539_),
    .A3(_08870_),
    .A4(_09687_),
    .ZN(_10540_));
 NAND4_X1 _20202_ (.A1(_10517_),
    .A2(_10525_),
    .A3(_10532_),
    .A4(_10540_),
    .ZN(_10541_));
 NOR2_X2 _20203_ (.A1(_10508_),
    .A2(_10541_),
    .ZN(_10542_));
 XNOR2_X1 _20204_ (.A(_10487_),
    .B(_10542_),
    .ZN(_10543_));
 XNOR2_X1 _20205_ (.A(_10543_),
    .B(_17094_),
    .ZN(_10544_));
 MUX2_X1 _20206_ (.A(_10311_),
    .B(_10544_),
    .S(_09040_),
    .Z(_00729_));
 XOR2_X1 _20207_ (.A(_17095_),
    .B(_17029_),
    .Z(_10545_));
 OAI21_X1 _20208_ (.A(_08646_),
    .B1(_08715_),
    .B2(_08698_),
    .ZN(_10546_));
 OAI211_X1 _20209_ (.A(_08523_),
    .B(_08615_),
    .C1(_09382_),
    .C2(_08794_),
    .ZN(_10547_));
 AND2_X1 _20210_ (.A1(_10546_),
    .A2(_10547_),
    .ZN(_10548_));
 OAI21_X1 _20211_ (.A(_08702_),
    .B1(_08681_),
    .B2(_09400_),
    .ZN(_10549_));
 AND4_X1 _20212_ (.A1(_08512_),
    .A2(_08506_),
    .A3(_08534_),
    .A4(_08675_),
    .ZN(_10550_));
 AOI211_X1 _20213_ (.A(_10550_),
    .B(_08738_),
    .C1(_08640_),
    .C2(_08513_),
    .ZN(_10551_));
 OAI21_X1 _20214_ (.A(_08702_),
    .B1(_08698_),
    .B2(_09810_),
    .ZN(_10552_));
 OAI21_X1 _20215_ (.A(_08513_),
    .B1(_08689_),
    .B2(_08758_),
    .ZN(_10553_));
 AND4_X1 _20216_ (.A1(_10549_),
    .A2(_10551_),
    .A3(_10552_),
    .A4(_10553_),
    .ZN(_10554_));
 OAI21_X1 _20217_ (.A(_08677_),
    .B1(_08685_),
    .B2(_08724_),
    .ZN(_10555_));
 OAI21_X1 _20218_ (.A(_08677_),
    .B1(_08732_),
    .B2(_08510_),
    .ZN(_10556_));
 AND4_X1 _20219_ (.A1(_10548_),
    .A2(_10554_),
    .A3(_10555_),
    .A4(_10556_),
    .ZN(_10557_));
 OAI21_X1 _20220_ (.A(_08650_),
    .B1(_08681_),
    .B2(_09400_),
    .ZN(_10558_));
 AOI21_X1 _20221_ (.A(_08754_),
    .B1(_08678_),
    .B2(_08557_),
    .ZN(_10559_));
 AOI21_X1 _20222_ (.A(_10559_),
    .B1(_08609_),
    .B2(_09543_),
    .ZN(_10560_));
 OAI211_X1 _20223_ (.A(_08609_),
    .B(_16706_),
    .C1(_08574_),
    .C2(_08515_),
    .ZN(_10561_));
 NOR2_X1 _20224_ (.A1(_09779_),
    .A2(_08756_),
    .ZN(_10562_));
 OAI21_X1 _20225_ (.A(_08572_),
    .B1(_08619_),
    .B2(_08606_),
    .ZN(_10563_));
 AND4_X1 _20226_ (.A1(_10560_),
    .A2(_10561_),
    .A3(_10562_),
    .A4(_10563_),
    .ZN(_10564_));
 AND2_X1 _20227_ (.A1(_08649_),
    .A2(_08575_),
    .ZN(_10565_));
 AND2_X1 _20228_ (.A1(_08649_),
    .A2(_08573_),
    .ZN(_10566_));
 AOI211_X1 _20229_ (.A(_10565_),
    .B(_10566_),
    .C1(_08650_),
    .C2(_09810_),
    .ZN(_10567_));
 AND2_X1 _20230_ (.A1(_08604_),
    .A2(_08578_),
    .ZN(_10568_));
 AOI21_X1 _20231_ (.A(_09572_),
    .B1(_09599_),
    .B2(_08680_),
    .ZN(_10569_));
 AOI211_X1 _20232_ (.A(_10568_),
    .B(_10569_),
    .C1(_08605_),
    .C2(_08732_),
    .ZN(_10570_));
 AND4_X1 _20233_ (.A1(_10558_),
    .A2(_10564_),
    .A3(_10567_),
    .A4(_10570_),
    .ZN(_10571_));
 OAI21_X1 _20234_ (.A(_08541_),
    .B1(_08621_),
    .B2(_08684_),
    .ZN(_10572_));
 OAI21_X1 _20235_ (.A(_08541_),
    .B1(_08527_),
    .B2(_08606_),
    .ZN(_10573_));
 OAI21_X1 _20236_ (.A(_08541_),
    .B1(_08679_),
    .B2(_08601_),
    .ZN(_10574_));
 AND3_X1 _20237_ (.A1(_10572_),
    .A2(_10573_),
    .A3(_10574_),
    .ZN(_10575_));
 AND2_X1 _20238_ (.A1(_08585_),
    .A2(_08575_),
    .ZN(_10576_));
 AND3_X1 _20239_ (.A1(_08688_),
    .A2(_08657_),
    .A3(_08581_),
    .ZN(_10577_));
 NOR4_X1 _20240_ (.A1(_10465_),
    .A2(_09536_),
    .A3(_10576_),
    .A4(_10577_),
    .ZN(_10578_));
 NAND2_X1 _20241_ (.A1(_09564_),
    .A2(_08622_),
    .ZN(_10579_));
 OAI21_X1 _20242_ (.A(_08622_),
    .B1(_08621_),
    .B2(_08684_),
    .ZN(_10580_));
 AND3_X1 _20243_ (.A1(_10579_),
    .A2(_10141_),
    .A3(_10580_),
    .ZN(_10581_));
 AND2_X1 _20244_ (.A1(_08573_),
    .A2(_08625_),
    .ZN(_10582_));
 AND2_X1 _20245_ (.A1(_08625_),
    .A2(_08640_),
    .ZN(_10583_));
 NOR4_X1 _20246_ (.A1(_10582_),
    .A2(_10467_),
    .A3(_10583_),
    .A4(_08627_),
    .ZN(_10584_));
 AND4_X1 _20247_ (.A1(_10575_),
    .A2(_10578_),
    .A3(_10581_),
    .A4(_10584_),
    .ZN(_10585_));
 AND2_X1 _20248_ (.A1(_08565_),
    .A2(_08553_),
    .ZN(_10586_));
 NAND3_X1 _20249_ (.A1(_08510_),
    .A2(_08632_),
    .A3(_08581_),
    .ZN(_10587_));
 NAND3_X1 _20250_ (.A1(_08640_),
    .A2(_08632_),
    .A3(_08563_),
    .ZN(_10588_));
 OAI211_X1 _20251_ (.A(_10587_),
    .B(_10588_),
    .C1(_08767_),
    .C2(_08802_),
    .ZN(_10589_));
 AND2_X1 _20252_ (.A1(_08564_),
    .A2(_08684_),
    .ZN(_10590_));
 OR4_X1 _20253_ (.A1(_10586_),
    .A2(_10589_),
    .A3(_10590_),
    .A4(_08772_),
    .ZN(_10591_));
 AND3_X1 _20254_ (.A1(_08588_),
    .A2(_08590_),
    .A3(_08629_),
    .ZN(_10592_));
 AND2_X1 _20255_ (.A1(_08697_),
    .A2(_08629_),
    .ZN(_10593_));
 AND4_X1 _20256_ (.A1(_08651_),
    .A2(_08631_),
    .A3(_08632_),
    .A4(_08512_),
    .ZN(_10594_));
 OR3_X1 _20257_ (.A1(_10592_),
    .A2(_10593_),
    .A3(_10594_),
    .ZN(_10595_));
 OAI21_X1 _20258_ (.A(_08664_),
    .B1(_08544_),
    .B2(_08665_),
    .ZN(_10596_));
 OAI211_X1 _20259_ (.A(_10596_),
    .B(_09818_),
    .C1(_09416_),
    .C2(_08802_),
    .ZN(_10597_));
 INV_X1 _20260_ (.A(_08765_),
    .ZN(_10598_));
 NAND2_X1 _20261_ (.A1(_08758_),
    .A2(_08549_),
    .ZN(_10599_));
 NAND3_X1 _20262_ (.A1(_08655_),
    .A2(_08642_),
    .A3(_08632_),
    .ZN(_10600_));
 NAND4_X1 _20263_ (.A1(_10598_),
    .A2(_08776_),
    .A3(_10599_),
    .A4(_10600_),
    .ZN(_10601_));
 NOR4_X1 _20264_ (.A1(_10591_),
    .A2(_10595_),
    .A3(_10597_),
    .A4(_10601_),
    .ZN(_10602_));
 NAND4_X1 _20265_ (.A1(_10557_),
    .A2(_10571_),
    .A3(_10585_),
    .A4(_10602_),
    .ZN(_10603_));
 NOR2_X2 _20266_ (.A1(_10603_),
    .A2(_08696_),
    .ZN(_10604_));
 OAI21_X1 _20267_ (.A(_08491_),
    .B1(_08454_),
    .B2(_10224_),
    .ZN(_10605_));
 AND3_X1 _20268_ (.A1(_08498_),
    .A2(_07992_),
    .A3(_07062_),
    .ZN(_10606_));
 OR3_X1 _20269_ (.A1(_09474_),
    .A2(_09466_),
    .A3(_10606_),
    .ZN(_10607_));
 OAI221_X1 _20270_ (.A(_10214_),
    .B1(_09304_),
    .B2(_09484_),
    .C1(_07641_),
    .C2(_07663_),
    .ZN(_10608_));
 AND2_X1 _20271_ (.A1(_08167_),
    .A2(_07828_),
    .ZN(_10609_));
 NAND2_X1 _20272_ (.A1(_10191_),
    .A2(_09906_),
    .ZN(_10610_));
 NOR4_X1 _20273_ (.A1(_10607_),
    .A2(_10608_),
    .A3(_10609_),
    .A4(_10610_),
    .ZN(_10611_));
 OAI21_X1 _20274_ (.A(_08491_),
    .B1(_09313_),
    .B2(_09837_),
    .ZN(_10612_));
 AOI21_X1 _20275_ (.A(_09311_),
    .B1(_09314_),
    .B2(_09838_),
    .ZN(_10613_));
 AOI211_X1 _20276_ (.A(_09524_),
    .B(_10613_),
    .C1(_07893_),
    .C2(_08337_),
    .ZN(_10614_));
 AND4_X1 _20277_ (.A1(_10605_),
    .A2(_10611_),
    .A3(_10612_),
    .A4(_10614_),
    .ZN(_10615_));
 AND2_X1 _20278_ (.A1(_07839_),
    .A2(_09289_),
    .ZN(_10616_));
 NOR4_X1 _20279_ (.A1(_09331_),
    .A2(_09357_),
    .A3(_07018_),
    .A4(_10616_),
    .ZN(_10617_));
 OR2_X1 _20280_ (.A1(_09321_),
    .A2(_07532_),
    .ZN(_10618_));
 OAI21_X1 _20281_ (.A(_07249_),
    .B1(_10618_),
    .B2(_09327_),
    .ZN(_10619_));
 OAI21_X1 _20282_ (.A(_08422_),
    .B1(_09321_),
    .B2(_08479_),
    .ZN(_10620_));
 OAI21_X1 _20283_ (.A(_07095_),
    .B1(_06952_),
    .B2(_07348_),
    .ZN(_10621_));
 AND3_X1 _20284_ (.A1(_10619_),
    .A2(_10620_),
    .A3(_10621_),
    .ZN(_10622_));
 OAI21_X1 _20285_ (.A(_07466_),
    .B1(_10224_),
    .B2(_09837_),
    .ZN(_10623_));
 OAI21_X1 _20286_ (.A(_09324_),
    .B1(_09352_),
    .B2(_08450_),
    .ZN(_10624_));
 AND4_X1 _20287_ (.A1(_09361_),
    .A2(_09868_),
    .A3(_10623_),
    .A4(_10624_),
    .ZN(_10625_));
 NAND4_X1 _20288_ (.A1(_10615_),
    .A2(_10617_),
    .A3(_10622_),
    .A4(_10625_),
    .ZN(_10626_));
 INV_X1 _20289_ (.A(_07040_),
    .ZN(_10627_));
 AOI21_X1 _20290_ (.A(_09468_),
    .B1(_08452_),
    .B2(_07707_),
    .ZN(_10628_));
 AOI21_X1 _20291_ (.A(_10628_),
    .B1(_07315_),
    .B2(_08337_),
    .ZN(_10629_));
 OAI211_X1 _20292_ (.A(_07315_),
    .B(_16714_),
    .C1(_08459_),
    .C2(_06908_),
    .ZN(_10630_));
 OAI21_X1 _20293_ (.A(_08014_),
    .B1(_08167_),
    .B2(_06952_),
    .ZN(_10631_));
 OAI21_X1 _20294_ (.A(_08014_),
    .B1(_07216_),
    .B2(_09456_),
    .ZN(_10632_));
 AND3_X1 _20295_ (.A1(_10631_),
    .A2(_10632_),
    .A3(_09854_),
    .ZN(_10633_));
 AND4_X1 _20296_ (.A1(_10627_),
    .A2(_10629_),
    .A3(_10630_),
    .A4(_10633_),
    .ZN(_10634_));
 AOI22_X1 _20297_ (.A1(_07029_),
    .A2(_09352_),
    .B1(_08156_),
    .B2(_08384_),
    .ZN(_10635_));
 AOI221_X1 _20298_ (.A(_09282_),
    .B1(_07948_),
    .B2(_07007_),
    .C1(_07348_),
    .C2(_07400_),
    .ZN(_10636_));
 AOI22_X1 _20299_ (.A1(_07095_),
    .A2(_09359_),
    .B1(_08413_),
    .B2(_08422_),
    .ZN(_10637_));
 AOI22_X1 _20300_ (.A1(_08485_),
    .A2(_07029_),
    .B1(_09327_),
    .B2(_08422_),
    .ZN(_10638_));
 AND4_X1 _20301_ (.A1(_10635_),
    .A2(_10636_),
    .A3(_10637_),
    .A4(_10638_),
    .ZN(_10639_));
 AOI21_X1 _20302_ (.A(_09277_),
    .B1(_09346_),
    .B2(_10373_),
    .ZN(_10640_));
 NOR4_X1 _20303_ (.A1(_10640_),
    .A2(_09504_),
    .A3(_09857_),
    .A4(_10375_),
    .ZN(_10641_));
 AOI22_X1 _20304_ (.A1(_08485_),
    .A2(_09456_),
    .B1(_07411_),
    .B2(_09272_),
    .ZN(_10642_));
 NAND2_X1 _20305_ (.A1(_08450_),
    .A2(_07904_),
    .ZN(_10643_));
 NAND3_X1 _20306_ (.A1(_07466_),
    .A2(_08384_),
    .A3(_09325_),
    .ZN(_10644_));
 NAND3_X1 _20307_ (.A1(_10642_),
    .A2(_10643_),
    .A3(_10644_),
    .ZN(_10645_));
 AOI21_X1 _20308_ (.A(_09261_),
    .B1(_08318_),
    .B2(_07510_),
    .ZN(_10646_));
 AOI21_X1 _20309_ (.A(_09261_),
    .B1(_09314_),
    .B2(_07970_),
    .ZN(_10647_));
 OAI21_X1 _20310_ (.A(_09525_),
    .B1(_07433_),
    .B2(_07488_),
    .ZN(_10648_));
 NOR4_X1 _20311_ (.A1(_10645_),
    .A2(_10646_),
    .A3(_10647_),
    .A4(_10648_),
    .ZN(_10649_));
 NAND4_X1 _20312_ (.A1(_10634_),
    .A2(_10639_),
    .A3(_10641_),
    .A4(_10649_),
    .ZN(_10650_));
 NOR2_X2 _20313_ (.A1(_10626_),
    .A2(_10650_),
    .ZN(_10651_));
 XOR2_X2 _20314_ (.A(_10604_),
    .B(_10651_),
    .Z(_10652_));
 OAI21_X1 _20315_ (.A(_09167_),
    .B1(_05114_),
    .B2(_04526_),
    .ZN(_10653_));
 AOI221_X4 _20316_ (.A(_10653_),
    .B1(_04888_),
    .B2(_05533_),
    .C1(_05907_),
    .C2(_04307_),
    .ZN(_10654_));
 OAI22_X1 _20317_ (.A1(_06215_),
    .A2(_09155_),
    .B1(_05114_),
    .B2(_05434_),
    .ZN(_10655_));
 AOI221_X4 _20318_ (.A(_10655_),
    .B1(_04636_),
    .B2(_05511_),
    .C1(_09612_),
    .C2(_05907_),
    .ZN(_10656_));
 AND2_X1 _20319_ (.A1(_05092_),
    .A2(_06556_),
    .ZN(_10657_));
 AOI221_X4 _20320_ (.A(_10657_),
    .B1(_06490_),
    .B2(_06391_),
    .C1(_04494_),
    .C2(_04307_),
    .ZN(_10658_));
 AND2_X1 _20321_ (.A1(_04263_),
    .A2(_09246_),
    .ZN(_10659_));
 NOR4_X1 _20322_ (.A1(_09192_),
    .A2(_09226_),
    .A3(_10659_),
    .A4(_10333_),
    .ZN(_10660_));
 AND4_X1 _20323_ (.A1(_10654_),
    .A2(_10656_),
    .A3(_10658_),
    .A4(_10660_),
    .ZN(_10661_));
 AOI22_X1 _20324_ (.A1(_06171_),
    .A2(_09615_),
    .B1(_05214_),
    .B2(_09612_),
    .ZN(_10662_));
 NOR4_X1 _20325_ (.A1(_09172_),
    .A2(_09173_),
    .A3(_09653_),
    .A4(_09216_),
    .ZN(_10663_));
 AND2_X1 _20326_ (.A1(_05907_),
    .A2(_04778_),
    .ZN(_10664_));
 NOR4_X1 _20327_ (.A1(_10355_),
    .A2(_10323_),
    .A3(_10664_),
    .A4(_10321_),
    .ZN(_10665_));
 AND4_X1 _20328_ (.A1(_05280_),
    .A2(_09643_),
    .A3(_10019_),
    .A4(_10022_),
    .ZN(_10666_));
 AND4_X1 _20329_ (.A1(_10662_),
    .A2(_10663_),
    .A3(_10665_),
    .A4(_10666_),
    .ZN(_10667_));
 OAI221_X1 _20330_ (.A(_05103_),
    .B1(_09197_),
    .B2(_05918_),
    .C1(_10016_),
    .C2(_06314_),
    .ZN(_10668_));
 AOI22_X1 _20331_ (.A1(_04614_),
    .A2(_10011_),
    .B1(_06446_),
    .B2(_09182_),
    .ZN(_10669_));
 OAI221_X1 _20332_ (.A(_10669_),
    .B1(_05203_),
    .B2(_10349_),
    .C1(_09185_),
    .C2(_04800_),
    .ZN(_10670_));
 NOR4_X1 _20333_ (.A1(_10668_),
    .A2(_09665_),
    .A3(_06666_),
    .A4(_10670_),
    .ZN(_10671_));
 NAND2_X1 _20334_ (.A1(_05045_),
    .A2(_04855_),
    .ZN(_10672_));
 NAND2_X1 _20335_ (.A1(_04494_),
    .A2(_06490_),
    .ZN(_10673_));
 AND4_X1 _20336_ (.A1(_10672_),
    .A2(_10328_),
    .A3(_09990_),
    .A4(_10673_),
    .ZN(_10674_));
 NAND2_X1 _20337_ (.A1(_05120_),
    .A2(_06446_),
    .ZN(_10675_));
 OAI21_X1 _20338_ (.A(_10675_),
    .B1(_04526_),
    .B2(_09238_),
    .ZN(_10676_));
 AND2_X1 _20339_ (.A1(_04559_),
    .A2(_05907_),
    .ZN(_10677_));
 NOR4_X1 _20340_ (.A1(_10676_),
    .A2(_10002_),
    .A3(_10677_),
    .A4(_09203_),
    .ZN(_10678_));
 NAND2_X1 _20341_ (.A1(_06160_),
    .A2(_05096_),
    .ZN(_10679_));
 NAND2_X1 _20342_ (.A1(_04844_),
    .A2(_04340_),
    .ZN(_10680_));
 AND4_X1 _20343_ (.A1(_09680_),
    .A2(_10679_),
    .A3(_10680_),
    .A4(_09625_),
    .ZN(_10681_));
 AOI22_X1 _20344_ (.A1(_04888_),
    .A2(_05599_),
    .B1(_04450_),
    .B2(_06556_),
    .ZN(_10682_));
 NAND2_X1 _20345_ (.A1(_04209_),
    .A2(_04778_),
    .ZN(_10683_));
 AND3_X1 _20346_ (.A1(_10682_),
    .A2(_10683_),
    .A3(_10075_),
    .ZN(_10684_));
 AND4_X1 _20347_ (.A1(_10674_),
    .A2(_10678_),
    .A3(_10681_),
    .A4(_10684_),
    .ZN(_10685_));
 NAND4_X1 _20348_ (.A1(_10661_),
    .A2(_10667_),
    .A3(_10671_),
    .A4(_10685_),
    .ZN(_10686_));
 NAND2_X1 _20349_ (.A1(_09178_),
    .A2(_09246_),
    .ZN(_10687_));
 AND2_X1 _20350_ (.A1(_05478_),
    .A2(_05775_),
    .ZN(_10688_));
 AOI221_X4 _20351_ (.A(_10688_),
    .B1(_05929_),
    .B2(_05511_),
    .C1(_06238_),
    .C2(_04614_),
    .ZN(_10689_));
 OAI21_X1 _20352_ (.A(_05522_),
    .B1(_09228_),
    .B2(_10011_),
    .ZN(_10690_));
 OAI21_X1 _20353_ (.A(_05786_),
    .B1(_05120_),
    .B2(_04340_),
    .ZN(_10691_));
 OAI21_X1 _20354_ (.A(_09246_),
    .B1(_06116_),
    .B2(_09623_),
    .ZN(_10692_));
 AND2_X1 _20355_ (.A1(_10691_),
    .A2(_10692_),
    .ZN(_10693_));
 AND4_X1 _20356_ (.A1(_10687_),
    .A2(_10689_),
    .A3(_10690_),
    .A4(_10693_),
    .ZN(_10694_));
 AND3_X1 _20357_ (.A1(_04767_),
    .A2(_04833_),
    .A3(_05110_),
    .ZN(_10695_));
 AND4_X1 _20358_ (.A1(_04950_),
    .A2(_05324_),
    .A3(_04329_),
    .A4(_04833_),
    .ZN(_10696_));
 AOI211_X1 _20359_ (.A(_10695_),
    .B(_10696_),
    .C1(_06238_),
    .C2(_05401_),
    .ZN(_10697_));
 AND2_X1 _20360_ (.A1(_05390_),
    .A2(_09182_),
    .ZN(_10698_));
 AOI211_X1 _20361_ (.A(_10698_),
    .B(_10316_),
    .C1(_05401_),
    .C2(_04537_),
    .ZN(_10699_));
 OAI21_X1 _20362_ (.A(_05632_),
    .B1(_09623_),
    .B2(_10011_),
    .ZN(_10700_));
 OAI211_X1 _20363_ (.A(_09158_),
    .B(_05874_),
    .C1(_05017_),
    .C2(_05445_),
    .ZN(_10701_));
 NAND4_X1 _20364_ (.A1(_09158_),
    .A2(_05203_),
    .A3(_06303_),
    .A4(_05874_),
    .ZN(_10702_));
 AND3_X1 _20365_ (.A1(_10700_),
    .A2(_10701_),
    .A3(_10702_),
    .ZN(_10703_));
 NAND4_X1 _20366_ (.A1(_10694_),
    .A2(_10697_),
    .A3(_10699_),
    .A4(_10703_),
    .ZN(_10704_));
 NOR2_X2 _20367_ (.A1(_10686_),
    .A2(_10704_),
    .ZN(_10705_));
 XNOR2_X1 _20368_ (.A(_10485_),
    .B(_10705_),
    .ZN(_10706_));
 XNOR2_X1 _20369_ (.A(_10652_),
    .B(_10706_),
    .ZN(_10707_));
 OR2_X1 _20370_ (.A1(_09102_),
    .A2(_09104_),
    .ZN(_10708_));
 INV_X1 _20371_ (.A(_10708_),
    .ZN(_10709_));
 AND3_X1 _20372_ (.A1(_08828_),
    .A2(_08874_),
    .A3(_08824_),
    .ZN(_10710_));
 AOI21_X1 _20373_ (.A(_10710_),
    .B1(_08829_),
    .B2(_09122_),
    .ZN(_10711_));
 NAND2_X1 _20374_ (.A1(_09004_),
    .A2(_09014_),
    .ZN(_10712_));
 NAND2_X1 _20375_ (.A1(_09025_),
    .A2(_08969_),
    .ZN(_10713_));
 NAND2_X1 _20376_ (.A1(_09046_),
    .A2(_09020_),
    .ZN(_10714_));
 AND4_X1 _20377_ (.A1(_10712_),
    .A2(_10713_),
    .A3(_09974_),
    .A4(_10714_),
    .ZN(_10715_));
 AND4_X1 _20378_ (.A1(_09024_),
    .A2(_10709_),
    .A3(_10711_),
    .A4(_10715_),
    .ZN(_10716_));
 AND4_X1 _20379_ (.A1(_09100_),
    .A2(_10716_),
    .A3(_09689_),
    .A4(_09693_),
    .ZN(_10717_));
 INV_X1 _20380_ (.A(_09074_),
    .ZN(_10718_));
 INV_X1 _20381_ (.A(_10251_),
    .ZN(_10719_));
 AOI21_X1 _20382_ (.A(_09143_),
    .B1(_10718_),
    .B2(_10719_),
    .ZN(_10720_));
 INV_X1 _20383_ (.A(_08941_),
    .ZN(_10721_));
 AOI21_X1 _20384_ (.A(_10721_),
    .B1(_10492_),
    .B2(_08991_),
    .ZN(_10722_));
 AND3_X1 _20385_ (.A1(_09026_),
    .A2(_08868_),
    .A3(_08867_),
    .ZN(_10723_));
 NOR4_X1 _20386_ (.A1(_10720_),
    .A2(_10722_),
    .A3(_09917_),
    .A4(_10723_),
    .ZN(_10724_));
 AND2_X1 _20387_ (.A1(_09106_),
    .A2(_08954_),
    .ZN(_10725_));
 AND2_X1 _20388_ (.A1(_09007_),
    .A2(_08965_),
    .ZN(_10726_));
 AND2_X1 _20389_ (.A1(_08911_),
    .A2(_08994_),
    .ZN(_10727_));
 AND3_X1 _20390_ (.A1(_08828_),
    .A2(_08964_),
    .A3(_08842_),
    .ZN(_10728_));
 NOR4_X1 _20391_ (.A1(_10725_),
    .A2(_10726_),
    .A3(_10727_),
    .A4(_10728_),
    .ZN(_10729_));
 AND2_X1 _20392_ (.A1(_08903_),
    .A2(_08994_),
    .ZN(_10730_));
 AND2_X1 _20393_ (.A1(_08838_),
    .A2(_08887_),
    .ZN(_10731_));
 NOR4_X1 _20394_ (.A1(_09140_),
    .A2(_10271_),
    .A3(_10730_),
    .A4(_10731_),
    .ZN(_10732_));
 AOI22_X1 _20395_ (.A1(_08982_),
    .A2(_09050_),
    .B1(_08969_),
    .B2(_08888_),
    .ZN(_10733_));
 AOI22_X1 _20396_ (.A1(_09031_),
    .A2(_08911_),
    .B1(_08847_),
    .B2(_09710_),
    .ZN(_10734_));
 AND4_X1 _20397_ (.A1(_10729_),
    .A2(_10732_),
    .A3(_10733_),
    .A4(_10734_),
    .ZN(_10735_));
 AND2_X1 _20398_ (.A1(_08906_),
    .A2(_09093_),
    .ZN(_10736_));
 AND2_X1 _20399_ (.A1(_08952_),
    .A2(_08915_),
    .ZN(_10737_));
 OR3_X1 _20400_ (.A1(_10736_),
    .A2(_10737_),
    .A3(_10501_),
    .ZN(_10738_));
 INV_X1 _20401_ (.A(_09752_),
    .ZN(_10739_));
 OAI21_X1 _20402_ (.A(_08865_),
    .B1(_09029_),
    .B2(_08894_),
    .ZN(_10740_));
 OAI211_X1 _20403_ (.A(_10739_),
    .B(_10740_),
    .C1(_09015_),
    .C2(_08932_),
    .ZN(_10741_));
 AOI21_X1 _20404_ (.A(_08932_),
    .B1(_08984_),
    .B2(_09061_),
    .ZN(_10742_));
 AOI21_X1 _20405_ (.A(_09109_),
    .B1(_09010_),
    .B2(_08875_),
    .ZN(_10743_));
 NOR4_X1 _20406_ (.A1(_10738_),
    .A2(_10741_),
    .A3(_10742_),
    .A4(_10743_),
    .ZN(_10744_));
 AND4_X1 _20407_ (.A1(_10717_),
    .A2(_10724_),
    .A3(_10735_),
    .A4(_10744_),
    .ZN(_10745_));
 AND2_X1 _20408_ (.A1(_09026_),
    .A2(_08909_),
    .ZN(_10746_));
 INV_X1 _20409_ (.A(_10746_),
    .ZN(_10747_));
 NAND2_X1 _20410_ (.A1(_08972_),
    .A2(_08989_),
    .ZN(_10748_));
 NAND2_X1 _20411_ (.A1(_09720_),
    .A2(_08987_),
    .ZN(_10749_));
 AOI22_X1 _20412_ (.A1(_09106_),
    .A2(_08945_),
    .B1(_08888_),
    .B2(_08909_),
    .ZN(_10750_));
 NAND4_X1 _20413_ (.A1(_10747_),
    .A2(_10748_),
    .A3(_10749_),
    .A4(_10750_),
    .ZN(_10751_));
 INV_X1 _20414_ (.A(_10276_),
    .ZN(_10752_));
 OAI21_X1 _20415_ (.A(_08982_),
    .B1(_09021_),
    .B2(_08969_),
    .ZN(_10753_));
 NAND2_X1 _20416_ (.A1(_10752_),
    .A2(_10753_),
    .ZN(_10754_));
 AOI21_X1 _20417_ (.A(_09057_),
    .B1(_10299_),
    .B2(_08984_),
    .ZN(_10755_));
 NOR4_X1 _20418_ (.A1(_10751_),
    .A2(_10754_),
    .A3(_09084_),
    .A4(_10755_),
    .ZN(_10756_));
 NAND2_X1 _20419_ (.A1(_09720_),
    .A2(_08943_),
    .ZN(_10757_));
 NAND4_X1 _20420_ (.A1(_08971_),
    .A2(_08959_),
    .A3(_10757_),
    .A4(_08955_),
    .ZN(_10758_));
 AOI21_X1 _20421_ (.A(_10758_),
    .B1(_08824_),
    .B2(_08839_),
    .ZN(_10759_));
 NAND2_X1 _20422_ (.A1(_09021_),
    .A2(_08829_),
    .ZN(_10760_));
 NAND2_X1 _20423_ (.A1(_08860_),
    .A2(_08829_),
    .ZN(_10761_));
 AND2_X1 _20424_ (.A1(_10760_),
    .A2(_10761_),
    .ZN(_10762_));
 NAND2_X1 _20425_ (.A1(_09720_),
    .A2(_08904_),
    .ZN(_10763_));
 OAI21_X1 _20426_ (.A(_09087_),
    .B1(_08998_),
    .B2(_08894_),
    .ZN(_10764_));
 AND4_X1 _20427_ (.A1(_08990_),
    .A2(_10762_),
    .A3(_10763_),
    .A4(_10764_),
    .ZN(_10765_));
 OR2_X1 _20428_ (.A1(_09072_),
    .A2(_09971_),
    .ZN(_10766_));
 AND2_X1 _20429_ (.A1(_09008_),
    .A2(_08998_),
    .ZN(_10767_));
 NOR4_X1 _20430_ (.A1(_10766_),
    .A2(_10302_),
    .A3(_09126_),
    .A4(_10767_),
    .ZN(_10768_));
 AND4_X1 _20431_ (.A1(_10756_),
    .A2(_10759_),
    .A3(_10765_),
    .A4(_10768_),
    .ZN(_10769_));
 NAND2_X2 _20432_ (.A1(_10745_),
    .A2(_10769_),
    .ZN(_10770_));
 XNOR2_X1 _20433_ (.A(_10707_),
    .B(_10770_),
    .ZN(_10771_));
 XNOR2_X1 _20434_ (.A(_10771_),
    .B(_17095_),
    .ZN(_10772_));
 MUX2_X1 _20435_ (.A(_10545_),
    .B(_10772_),
    .S(_09040_),
    .Z(_00730_));
 AND2_X1 _20436_ (.A1(_07400_),
    .A2(_09272_),
    .ZN(_10773_));
 AOI21_X1 _20437_ (.A(_10373_),
    .B1(_09287_),
    .B2(_10385_),
    .ZN(_10774_));
 AOI211_X1 _20438_ (.A(_10773_),
    .B(_10774_),
    .C1(_08498_),
    .C2(_07400_),
    .ZN(_10775_));
 NAND2_X1 _20439_ (.A1(_09887_),
    .A2(_08014_),
    .ZN(_10776_));
 OAI21_X1 _20440_ (.A(_08014_),
    .B1(_07762_),
    .B2(_07904_),
    .ZN(_10777_));
 OAI21_X1 _20441_ (.A(_08014_),
    .B1(_09330_),
    .B2(_09288_),
    .ZN(_10778_));
 OAI211_X1 _20442_ (.A(_08189_),
    .B(_08463_),
    .C1(_07609_),
    .C2(_07378_),
    .ZN(_10779_));
 AND4_X1 _20443_ (.A1(_10776_),
    .A2(_10777_),
    .A3(_10778_),
    .A4(_10779_),
    .ZN(_10780_));
 OAI21_X1 _20444_ (.A(_06732_),
    .B1(_09887_),
    .B2(_07751_),
    .ZN(_10781_));
 AND2_X1 _20445_ (.A1(_07861_),
    .A2(_07828_),
    .ZN(_10782_));
 AND2_X1 _20446_ (.A1(_07828_),
    .A2(_07872_),
    .ZN(_10783_));
 NOR4_X1 _20447_ (.A1(_10782_),
    .A2(_10609_),
    .A3(_09856_),
    .A4(_10783_),
    .ZN(_10784_));
 NAND4_X1 _20448_ (.A1(_10775_),
    .A2(_10780_),
    .A3(_10781_),
    .A4(_10784_),
    .ZN(_10785_));
 AND3_X1 _20449_ (.A1(_07674_),
    .A2(_08458_),
    .A3(_07183_),
    .ZN(_10786_));
 OR4_X1 _20450_ (.A1(_09338_),
    .A2(_10199_),
    .A3(_10786_),
    .A4(_09339_),
    .ZN(_10787_));
 OAI21_X1 _20451_ (.A(_07084_),
    .B1(_07216_),
    .B2(_09456_),
    .ZN(_10788_));
 OAI21_X1 _20452_ (.A(_07084_),
    .B1(_07904_),
    .B2(_06776_),
    .ZN(_10789_));
 NAND3_X1 _20453_ (.A1(_10788_),
    .A2(_10789_),
    .A3(_09507_),
    .ZN(_10790_));
 OAI21_X1 _20454_ (.A(_08145_),
    .B1(_08308_),
    .B2(_07784_),
    .ZN(_10791_));
 NAND4_X1 _20455_ (.A1(_08189_),
    .A2(_07062_),
    .A3(_08091_),
    .A4(_08478_),
    .ZN(_10792_));
 AND2_X1 _20456_ (.A1(_10791_),
    .A2(_10792_),
    .ZN(_10793_));
 OAI21_X1 _20457_ (.A(_08145_),
    .B1(_09348_),
    .B2(_07609_),
    .ZN(_10794_));
 OAI21_X1 _20458_ (.A(_07893_),
    .B1(_09321_),
    .B2(_07532_),
    .ZN(_10795_));
 OAI21_X1 _20459_ (.A(_07893_),
    .B1(_09289_),
    .B2(_08455_),
    .ZN(_10796_));
 NAND4_X1 _20460_ (.A1(_10793_),
    .A2(_10794_),
    .A3(_10795_),
    .A4(_10796_),
    .ZN(_10797_));
 NOR4_X1 _20461_ (.A1(_10785_),
    .A2(_10787_),
    .A3(_10790_),
    .A4(_10797_),
    .ZN(_10798_));
 AOI211_X1 _20462_ (.A(_06842_),
    .B(_07293_),
    .C1(_06754_),
    .C2(_08091_),
    .ZN(_10799_));
 OAI21_X1 _20463_ (.A(_07565_),
    .B1(_06952_),
    .B2(_07872_),
    .ZN(_10800_));
 OAI211_X1 _20464_ (.A(_10800_),
    .B(_09892_),
    .C1(_09261_),
    .C2(_10385_),
    .ZN(_10801_));
 NAND4_X1 _20465_ (.A1(_08069_),
    .A2(_06974_),
    .A3(_07543_),
    .A4(_08403_),
    .ZN(_10802_));
 OAI211_X1 _20466_ (.A(_09268_),
    .B(_10802_),
    .C1(_09287_),
    .C2(_07293_),
    .ZN(_10803_));
 AND2_X1 _20467_ (.A1(_07850_),
    .A2(_06919_),
    .ZN(_10804_));
 AND2_X1 _20468_ (.A1(_10804_),
    .A2(_07007_),
    .ZN(_10805_));
 NOR4_X1 _20469_ (.A1(_10799_),
    .A2(_10801_),
    .A3(_10803_),
    .A4(_10805_),
    .ZN(_10806_));
 AOI221_X4 _20470_ (.A(_07641_),
    .B1(_06754_),
    .B2(_08458_),
    .C1(_07128_),
    .C2(_07740_),
    .ZN(_10807_));
 AND2_X1 _20471_ (.A1(_06831_),
    .A2(_07696_),
    .ZN(_10808_));
 OR2_X1 _20472_ (.A1(_08471_),
    .A2(_10808_),
    .ZN(_10809_));
 NOR2_X1 _20473_ (.A1(_08047_),
    .A2(_09289_),
    .ZN(_10810_));
 NOR2_X1 _20474_ (.A1(_10810_),
    .A2(_09468_),
    .ZN(_10811_));
 AND2_X1 _20475_ (.A1(_07631_),
    .A2(_07029_),
    .ZN(_10812_));
 NOR4_X1 _20476_ (.A1(_10807_),
    .A2(_10809_),
    .A3(_10811_),
    .A4(_10812_),
    .ZN(_10813_));
 INV_X1 _20477_ (.A(_10221_),
    .ZN(_10814_));
 AND3_X1 _20478_ (.A1(_09490_),
    .A2(_09906_),
    .A3(_09284_),
    .ZN(_10815_));
 OAI21_X1 _20479_ (.A(_07238_),
    .B1(_10804_),
    .B2(_07029_),
    .ZN(_10816_));
 OAI21_X1 _20480_ (.A(_08490_),
    .B1(_09324_),
    .B2(_07948_),
    .ZN(_10817_));
 AND4_X1 _20481_ (.A1(_10814_),
    .A2(_10815_),
    .A3(_10816_),
    .A4(_10817_),
    .ZN(_10818_));
 OAI21_X1 _20482_ (.A(_09352_),
    .B1(_10404_),
    .B2(_09348_),
    .ZN(_10819_));
 OAI21_X1 _20483_ (.A(_07466_),
    .B1(_08454_),
    .B2(_08308_),
    .ZN(_10820_));
 OAI211_X1 _20484_ (.A(_08189_),
    .B(_08211_),
    .C1(_08167_),
    .C2(_09272_),
    .ZN(_10821_));
 AND4_X1 _20485_ (.A1(_09463_),
    .A2(_10819_),
    .A3(_10820_),
    .A4(_10821_),
    .ZN(_10822_));
 AND4_X1 _20486_ (.A1(_10806_),
    .A2(_10813_),
    .A3(_10818_),
    .A4(_10822_),
    .ZN(_10823_));
 AND2_X2 _20487_ (.A1(_10798_),
    .A2(_10823_),
    .ZN(_10824_));
 NAND2_X1 _20488_ (.A1(_04537_),
    .A2(_05522_),
    .ZN(_10825_));
 AOI21_X1 _20489_ (.A(_05114_),
    .B1(_09200_),
    .B2(_09201_),
    .ZN(_10826_));
 NOR2_X1 _20490_ (.A1(_10056_),
    .A2(_10826_),
    .ZN(_10827_));
 OAI21_X1 _20491_ (.A(_05214_),
    .B1(_05064_),
    .B2(_04450_),
    .ZN(_10828_));
 OAI21_X1 _20492_ (.A(_05522_),
    .B1(_05929_),
    .B2(_09178_),
    .ZN(_10829_));
 AND4_X1 _20493_ (.A1(_10825_),
    .A2(_10827_),
    .A3(_10828_),
    .A4(_10829_),
    .ZN(_10830_));
 OAI21_X1 _20494_ (.A(_09246_),
    .B1(_09615_),
    .B2(_10008_),
    .ZN(_10831_));
 OAI21_X1 _20495_ (.A(_05896_),
    .B1(_05676_),
    .B2(_04778_),
    .ZN(_10832_));
 NAND2_X1 _20496_ (.A1(_09178_),
    .A2(_05896_),
    .ZN(_10833_));
 AND3_X1 _20497_ (.A1(_10832_),
    .A2(_10833_),
    .A3(_09605_),
    .ZN(_10834_));
 OAI21_X1 _20498_ (.A(_09246_),
    .B1(_04307_),
    .B2(_06413_),
    .ZN(_10835_));
 OAI221_X1 _20499_ (.A(_05907_),
    .B1(_05137_),
    .B2(_05192_),
    .C1(_09612_),
    .C2(_05863_),
    .ZN(_10836_));
 AND4_X1 _20500_ (.A1(_10831_),
    .A2(_10834_),
    .A3(_10835_),
    .A4(_10836_),
    .ZN(_10837_));
 OAI211_X1 _20501_ (.A(_09158_),
    .B(_05874_),
    .C1(_05096_),
    .C2(_04636_),
    .ZN(_10838_));
 NAND4_X1 _20502_ (.A1(_10366_),
    .A2(_10107_),
    .A3(_05643_),
    .A4(_10838_),
    .ZN(_10839_));
 NOR2_X1 _20503_ (.A1(_09238_),
    .A2(_04526_),
    .ZN(_10840_));
 NAND3_X1 _20504_ (.A1(_05775_),
    .A2(_04713_),
    .A3(_05313_),
    .ZN(_10841_));
 OAI211_X1 _20505_ (.A(_10841_),
    .B(_09628_),
    .C1(_05456_),
    .C2(_09238_),
    .ZN(_10842_));
 AOI21_X1 _20506_ (.A(_09238_),
    .B1(_09185_),
    .B2(_05170_),
    .ZN(_10843_));
 NOR4_X1 _20507_ (.A1(_10839_),
    .A2(_10840_),
    .A3(_10842_),
    .A4(_10843_),
    .ZN(_10844_));
 NOR4_X1 _20508_ (.A1(_05412_),
    .A2(_09151_),
    .A3(_10698_),
    .A4(_10695_),
    .ZN(_10845_));
 OAI221_X1 _20509_ (.A(_05291_),
    .B1(_04959_),
    .B2(_05192_),
    .C1(_05863_),
    .C2(_05797_),
    .ZN(_10846_));
 AND3_X1 _20510_ (.A1(_10845_),
    .A2(_10324_),
    .A3(_10846_),
    .ZN(_10847_));
 NAND4_X2 _20511_ (.A1(_10830_),
    .A2(_10837_),
    .A3(_10844_),
    .A4(_10847_),
    .ZN(_10848_));
 NAND2_X1 _20512_ (.A1(_06160_),
    .A2(_04537_),
    .ZN(_10849_));
 NAND4_X1 _20513_ (.A1(_09225_),
    .A2(_09651_),
    .A3(_10849_),
    .A4(_10679_),
    .ZN(_10850_));
 AOI211_X1 _20514_ (.A(_06402_),
    .B(_06215_),
    .C1(_05137_),
    .C2(_04680_),
    .ZN(_10851_));
 NOR2_X1 _20515_ (.A1(_10075_),
    .A2(_05313_),
    .ZN(_10852_));
 OAI21_X1 _20516_ (.A(_06270_),
    .B1(_04340_),
    .B2(_04746_),
    .ZN(_10853_));
 NAND3_X1 _20517_ (.A1(_10853_),
    .A2(_09996_),
    .A3(_09995_),
    .ZN(_10854_));
 NOR4_X1 _20518_ (.A1(_10850_),
    .A2(_10851_),
    .A3(_10852_),
    .A4(_10854_),
    .ZN(_10855_));
 OAI21_X1 _20519_ (.A(_04209_),
    .B1(_09615_),
    .B2(_05159_),
    .ZN(_10856_));
 NAND4_X1 _20520_ (.A1(_10856_),
    .A2(_10349_),
    .A3(_10683_),
    .A4(_04351_),
    .ZN(_10857_));
 OAI211_X1 _20521_ (.A(_10088_),
    .B(_10680_),
    .C1(_09193_),
    .C2(_09189_),
    .ZN(_10858_));
 NOR4_X1 _20522_ (.A1(_10857_),
    .A2(_10858_),
    .A3(_09192_),
    .A4(_10086_),
    .ZN(_10859_));
 AOI21_X1 _20523_ (.A(_09197_),
    .B1(_09170_),
    .B2(_09201_),
    .ZN(_10860_));
 OAI211_X1 _20524_ (.A(_10093_),
    .B(_10344_),
    .C1(_09197_),
    .C2(_09189_),
    .ZN(_10861_));
 AOI21_X1 _20525_ (.A(_04800_),
    .B1(_05126_),
    .B2(_09198_),
    .ZN(_10862_));
 AOI21_X1 _20526_ (.A(_04800_),
    .B1(_09183_),
    .B2(_09608_),
    .ZN(_10863_));
 NOR4_X1 _20527_ (.A1(_10860_),
    .A2(_10861_),
    .A3(_10862_),
    .A4(_10863_),
    .ZN(_10864_));
 OAI21_X1 _20528_ (.A(_06556_),
    .B1(_09182_),
    .B2(_10008_),
    .ZN(_10865_));
 OAI21_X1 _20529_ (.A(_06446_),
    .B1(_06468_),
    .B2(_09623_),
    .ZN(_10866_));
 OAI21_X1 _20530_ (.A(_06391_),
    .B1(_05064_),
    .B2(_06413_),
    .ZN(_10867_));
 OAI211_X1 _20531_ (.A(_06556_),
    .B(_04680_),
    .C1(_06303_),
    .C2(_04950_),
    .ZN(_10868_));
 AND4_X1 _20532_ (.A1(_10865_),
    .A2(_10866_),
    .A3(_10867_),
    .A4(_10868_),
    .ZN(_10869_));
 NAND4_X2 _20533_ (.A1(_10855_),
    .A2(_10859_),
    .A3(_10864_),
    .A4(_10869_),
    .ZN(_10870_));
 NOR2_X4 _20534_ (.A1(_10848_),
    .A2(_10870_),
    .ZN(_10871_));
 XOR2_X2 _20535_ (.A(_10824_),
    .B(_10871_),
    .Z(_10872_));
 OAI21_X1 _20536_ (.A(_09031_),
    .B1(_09014_),
    .B2(_08989_),
    .ZN(_10873_));
 OAI21_X1 _20537_ (.A(_10873_),
    .B1(_10718_),
    .B2(_09097_),
    .ZN(_10874_));
 OR4_X1 _20538_ (.A1(_09023_),
    .A2(_10874_),
    .A3(_10276_),
    .A4(_09977_),
    .ZN(_10875_));
 AND2_X1 _20539_ (.A1(_10303_),
    .A2(_09116_),
    .ZN(_10876_));
 OR4_X1 _20540_ (.A1(_09958_),
    .A2(_10876_),
    .A3(_09959_),
    .A4(_10726_),
    .ZN(_10877_));
 OAI21_X1 _20541_ (.A(_09005_),
    .B1(_09017_),
    .B2(_09690_),
    .ZN(_10878_));
 OAI21_X1 _20542_ (.A(_09005_),
    .B1(_08860_),
    .B2(_08855_),
    .ZN(_10879_));
 OAI211_X1 _20543_ (.A(_10878_),
    .B(_10879_),
    .C1(_09109_),
    .C2(_10719_),
    .ZN(_10880_));
 OR4_X1 _20544_ (.A1(_09027_),
    .A2(_10270_),
    .A3(_10746_),
    .A4(_09740_),
    .ZN(_10881_));
 NOR4_X1 _20545_ (.A1(_10875_),
    .A2(_10877_),
    .A3(_10880_),
    .A4(_10881_),
    .ZN(_10882_));
 AND3_X1 _20546_ (.A1(_08882_),
    .A2(_08827_),
    .A3(_08914_),
    .ZN(_10883_));
 AND3_X1 _20547_ (.A1(_09062_),
    .A2(_08873_),
    .A3(_08941_),
    .ZN(_10884_));
 AOI211_X1 _20548_ (.A(_10883_),
    .B(_10884_),
    .C1(_10251_),
    .C2(_08941_),
    .ZN(_10885_));
 NAND2_X1 _20549_ (.A1(_08936_),
    .A2(_09077_),
    .ZN(_10886_));
 AND4_X1 _20550_ (.A1(_10886_),
    .A2(_10257_),
    .A3(_09117_),
    .A4(_09737_),
    .ZN(_10887_));
 NAND2_X1 _20551_ (.A1(_09106_),
    .A2(_08998_),
    .ZN(_10888_));
 OAI211_X1 _20552_ (.A(_08913_),
    .B(_08914_),
    .C1(_09710_),
    .C2(_08989_),
    .ZN(_10889_));
 NAND2_X1 _20553_ (.A1(_09106_),
    .A2(_09009_),
    .ZN(_10890_));
 AND4_X1 _20554_ (.A1(_10888_),
    .A2(_10889_),
    .A3(_10890_),
    .A4(_09119_),
    .ZN(_10891_));
 AND2_X1 _20555_ (.A1(_08901_),
    .A2(_08903_),
    .ZN(_10892_));
 INV_X1 _20556_ (.A(_10892_),
    .ZN(_10893_));
 NAND3_X1 _20557_ (.A1(_09048_),
    .A2(_08886_),
    .A3(_08914_),
    .ZN(_10894_));
 AND4_X1 _20558_ (.A1(_10893_),
    .A2(_08921_),
    .A3(_08925_),
    .A4(_10894_),
    .ZN(_10895_));
 AND4_X1 _20559_ (.A1(_10885_),
    .A2(_10887_),
    .A3(_10891_),
    .A4(_10895_),
    .ZN(_10896_));
 OAI21_X1 _20560_ (.A(_08830_),
    .B1(_08986_),
    .B2(_09050_),
    .ZN(_10897_));
 AND4_X1 _20561_ (.A1(_10528_),
    .A2(_09944_),
    .A3(_09938_),
    .A4(_10897_),
    .ZN(_10898_));
 NAND2_X1 _20562_ (.A1(_08907_),
    .A2(_08847_),
    .ZN(_10899_));
 AND3_X1 _20563_ (.A1(_10899_),
    .A2(_09703_),
    .A3(_08861_),
    .ZN(_10900_));
 OAI211_X1 _20564_ (.A(_08847_),
    .B(_09107_),
    .C1(_09115_),
    .C2(_08858_),
    .ZN(_10901_));
 AND4_X1 _20565_ (.A1(_10241_),
    .A2(_10900_),
    .A3(_10243_),
    .A4(_10901_),
    .ZN(_10902_));
 NAND2_X1 _20566_ (.A1(_09075_),
    .A2(_08853_),
    .ZN(_10903_));
 NAND2_X1 _20567_ (.A1(_09075_),
    .A2(_08943_),
    .ZN(_10904_));
 AND4_X1 _20568_ (.A1(_08881_),
    .A2(_10534_),
    .A3(_10903_),
    .A4(_10904_),
    .ZN(_10905_));
 NAND2_X1 _20569_ (.A1(_10266_),
    .A2(_09138_),
    .ZN(_10906_));
 AOI211_X1 _20570_ (.A(_08890_),
    .B(_10906_),
    .C1(_08888_),
    .C2(_08969_),
    .ZN(_10907_));
 AND4_X1 _20571_ (.A1(_10898_),
    .A2(_10902_),
    .A3(_10905_),
    .A4(_10907_),
    .ZN(_10908_));
 OAI21_X1 _20572_ (.A(_09053_),
    .B1(_08911_),
    .B2(_08943_),
    .ZN(_10909_));
 INV_X1 _20573_ (.A(_09748_),
    .ZN(_10910_));
 NAND2_X1 _20574_ (.A1(_08903_),
    .A2(_09053_),
    .ZN(_10911_));
 AND3_X1 _20575_ (.A1(_10910_),
    .A2(_08960_),
    .A3(_10911_),
    .ZN(_10912_));
 AND4_X1 _20576_ (.A1(_08822_),
    .A2(_08833_),
    .A3(_09107_),
    .A4(_08950_),
    .ZN(_10913_));
 AOI21_X1 _20577_ (.A(_10913_),
    .B1(_09017_),
    .B2(_08972_),
    .ZN(_10914_));
 OAI21_X1 _20578_ (.A(_08972_),
    .B1(_08882_),
    .B2(_10251_),
    .ZN(_10915_));
 AND4_X1 _20579_ (.A1(_10909_),
    .A2(_10912_),
    .A3(_10914_),
    .A4(_10915_),
    .ZN(_10916_));
 OAI21_X1 _20580_ (.A(_08982_),
    .B1(_08998_),
    .B2(_08989_),
    .ZN(_10917_));
 NOR3_X1 _20581_ (.A1(_09951_),
    .A2(_08978_),
    .A3(_09044_),
    .ZN(_10918_));
 OAI21_X1 _20582_ (.A(_09087_),
    .B1(_08882_),
    .B2(_09046_),
    .ZN(_10919_));
 OAI211_X1 _20583_ (.A(_09087_),
    .B(_09107_),
    .C1(_08973_),
    .C2(_08878_),
    .ZN(_10920_));
 AND2_X1 _20584_ (.A1(_10919_),
    .A2(_10920_),
    .ZN(_10921_));
 AND4_X1 _20585_ (.A1(_10916_),
    .A2(_10917_),
    .A3(_10918_),
    .A4(_10921_),
    .ZN(_10922_));
 NAND4_X1 _20586_ (.A1(_10882_),
    .A2(_10896_),
    .A3(_10908_),
    .A4(_10922_),
    .ZN(_10923_));
 NOR2_X2 _20587_ (.A1(_10923_),
    .A2(_09752_),
    .ZN(_10924_));
 XOR2_X1 _20588_ (.A(_10872_),
    .B(_10924_),
    .Z(_10925_));
 XNOR2_X1 _20589_ (.A(_10604_),
    .B(_08811_),
    .ZN(_10926_));
 OAI21_X1 _20590_ (.A(_09038_),
    .B1(_10925_),
    .B2(_10926_),
    .ZN(_10927_));
 AOI21_X1 _20591_ (.A(_10927_),
    .B1(_10926_),
    .B2(_10925_),
    .ZN(_10928_));
 AND2_X1 _20592_ (.A1(_01331_),
    .A2(_17040_),
    .ZN(_10929_));
 NOR2_X1 _20593_ (.A1(_10928_),
    .A2(_10929_),
    .ZN(_10930_));
 XNOR2_X1 _20594_ (.A(_10930_),
    .B(_17096_),
    .ZN(_00731_));
 CLKBUF_X2 _20595_ (.A(_17097_),
    .Z(_10931_));
 BUF_X2 _20596_ (.A(_10931_),
    .Z(_10932_));
 XOR2_X1 _20597_ (.A(_17051_),
    .B(_10932_),
    .Z(_10933_));
 XNOR2_X1 _20598_ (.A(_08502_),
    .B(_08722_),
    .ZN(_10934_));
 XOR2_X1 _20599_ (.A(_10871_),
    .B(_01049_),
    .Z(_10935_));
 XNOR2_X1 _20600_ (.A(_10934_),
    .B(_10935_),
    .ZN(_10936_));
 XOR2_X1 _20601_ (.A(_10936_),
    .B(_09148_),
    .Z(_10937_));
 MUX2_X1 _20602_ (.A(_10933_),
    .B(_10937_),
    .S(_09040_),
    .Z(_00692_));
 BUF_X2 _20603_ (.A(_17098_),
    .Z(_10938_));
 XOR2_X1 _20604_ (.A(_10938_),
    .B(_17062_),
    .Z(_10939_));
 XNOR2_X1 _20605_ (.A(_09148_),
    .B(_09759_),
    .ZN(_10940_));
 XOR2_X2 _20606_ (.A(_06677_),
    .B(_10871_),
    .Z(_10941_));
 XNOR2_X1 _20607_ (.A(_10941_),
    .B(_09448_),
    .ZN(_10942_));
 XNOR2_X1 _20608_ (.A(_10940_),
    .B(_10942_),
    .ZN(_10943_));
 INV_X1 _20609_ (.A(_17098_),
    .ZN(_10944_));
 CLKBUF_X2 _20610_ (.A(_10944_),
    .Z(_10945_));
 BUF_X2 _20611_ (.A(_10945_),
    .Z(_10946_));
 XNOR2_X1 _20612_ (.A(_10943_),
    .B(_10946_),
    .ZN(_10947_));
 MUX2_X1 _20613_ (.A(_10939_),
    .B(_10947_),
    .S(_09040_),
    .Z(_00693_));
 XOR2_X1 _20614_ (.A(_17068_),
    .B(_16946_),
    .Z(_10948_));
 XNOR2_X1 _20615_ (.A(_09258_),
    .B(_09758_),
    .ZN(_10949_));
 XOR2_X1 _20616_ (.A(_09604_),
    .B(_10949_),
    .Z(_10950_));
 XNOR2_X1 _20617_ (.A(_10950_),
    .B(_09984_),
    .ZN(_10951_));
 XNOR2_X1 _20618_ (.A(_10951_),
    .B(_17068_),
    .ZN(_10952_));
 MUX2_X1 _20619_ (.A(_10948_),
    .B(_10952_),
    .S(_09040_),
    .Z(_00694_));
 XOR2_X1 _20620_ (.A(_17069_),
    .B(_16957_),
    .Z(_10953_));
 XNOR2_X1 _20621_ (.A(_09685_),
    .B(_10871_),
    .ZN(_10954_));
 XNOR2_X1 _20622_ (.A(_10954_),
    .B(_10307_),
    .ZN(_10955_));
 XNOR2_X1 _20623_ (.A(_09986_),
    .B(_10955_),
    .ZN(_10956_));
 XNOR2_X1 _20624_ (.A(_10956_),
    .B(_17069_),
    .ZN(_10957_));
 BUF_X2 _20625_ (.A(_09039_),
    .Z(_10958_));
 MUX2_X1 _20626_ (.A(_10953_),
    .B(_10957_),
    .S(_10958_),
    .Z(_00695_));
 XOR2_X1 _20627_ (.A(_17070_),
    .B(_16966_),
    .Z(_10959_));
 XOR2_X2 _20628_ (.A(_10060_),
    .B(_10871_),
    .Z(_10960_));
 XNOR2_X1 _20629_ (.A(_10960_),
    .B(_10238_),
    .ZN(_10961_));
 XNOR2_X1 _20630_ (.A(_10308_),
    .B(_10542_),
    .ZN(_10962_));
 XNOR2_X1 _20631_ (.A(_10961_),
    .B(_10962_),
    .ZN(_10963_));
 INV_X1 _20632_ (.A(_17070_),
    .ZN(_10964_));
 XNOR2_X1 _20633_ (.A(_10963_),
    .B(_10964_),
    .ZN(_10965_));
 MUX2_X1 _20634_ (.A(_10959_),
    .B(_10965_),
    .S(_10958_),
    .Z(_00696_));
 XOR2_X1 _20635_ (.A(_17071_),
    .B(_16967_),
    .Z(_10966_));
 XNOR2_X1 _20636_ (.A(_10542_),
    .B(_10119_),
    .ZN(_10967_));
 XNOR2_X1 _20637_ (.A(_10967_),
    .B(_10770_),
    .ZN(_10968_));
 XNOR2_X1 _20638_ (.A(_10968_),
    .B(_10486_),
    .ZN(_10969_));
 INV_X1 _20639_ (.A(_17071_),
    .ZN(_10970_));
 XNOR2_X1 _20640_ (.A(_10969_),
    .B(_10970_),
    .ZN(_10971_));
 MUX2_X1 _20641_ (.A(_10966_),
    .B(_10971_),
    .S(_10958_),
    .Z(_00697_));
 XOR2_X1 _20642_ (.A(_17072_),
    .B(_16968_),
    .Z(_10972_));
 XOR2_X1 _20643_ (.A(_10770_),
    .B(_10371_),
    .Z(_10973_));
 XNOR2_X1 _20644_ (.A(_10973_),
    .B(_10652_),
    .ZN(_10974_));
 XNOR2_X1 _20645_ (.A(_10974_),
    .B(_10924_),
    .ZN(_10975_));
 INV_X1 _20646_ (.A(_17072_),
    .ZN(_10976_));
 XNOR2_X1 _20647_ (.A(_10975_),
    .B(_10976_),
    .ZN(_10977_));
 MUX2_X1 _20648_ (.A(_10972_),
    .B(_10977_),
    .S(_10958_),
    .Z(_00698_));
 XOR2_X1 _20649_ (.A(_17073_),
    .B(_16969_),
    .Z(_10978_));
 XNOR2_X1 _20650_ (.A(_10705_),
    .B(_08811_),
    .ZN(_10979_));
 INV_X1 _20651_ (.A(_10824_),
    .ZN(_10980_));
 XNOR2_X1 _20652_ (.A(_10979_),
    .B(_10980_),
    .ZN(_10981_));
 XNOR2_X1 _20653_ (.A(_10924_),
    .B(_09035_),
    .ZN(_10982_));
 XNOR2_X1 _20654_ (.A(_10981_),
    .B(_10982_),
    .ZN(_10983_));
 INV_X1 _20655_ (.A(_17073_),
    .ZN(_10984_));
 XNOR2_X1 _20656_ (.A(_10983_),
    .B(_10984_),
    .ZN(_10985_));
 MUX2_X1 _20657_ (.A(_10978_),
    .B(_10985_),
    .S(_10958_),
    .Z(_00699_));
 CLKBUF_X2 _20658_ (.A(_17074_),
    .Z(_10986_));
 BUF_X2 _20659_ (.A(_10986_),
    .Z(_10987_));
 XOR2_X1 _20660_ (.A(_16970_),
    .B(_10987_),
    .Z(_10988_));
 XNOR2_X1 _20661_ (.A(_06677_),
    .B(_01050_),
    .ZN(_10989_));
 XNOR2_X1 _20662_ (.A(_10989_),
    .B(_10872_),
    .ZN(_10990_));
 XNOR2_X1 _20663_ (.A(_09147_),
    .B(_08722_),
    .ZN(_10991_));
 XNOR2_X1 _20664_ (.A(_10990_),
    .B(_10991_),
    .ZN(_10992_));
 MUX2_X1 _20665_ (.A(_10988_),
    .B(_10992_),
    .S(_10958_),
    .Z(_00660_));
 BUF_X2 _20666_ (.A(_17075_),
    .Z(_10993_));
 XOR2_X1 _20667_ (.A(_16971_),
    .B(_10993_),
    .Z(_10994_));
 XNOR2_X1 _20668_ (.A(_10941_),
    .B(_10949_),
    .ZN(_10995_));
 XNOR2_X1 _20669_ (.A(_09447_),
    .B(_01051_),
    .ZN(_10996_));
 XNOR2_X2 _20670_ (.A(_08502_),
    .B(_10824_),
    .ZN(_10997_));
 XNOR2_X1 _20671_ (.A(_10996_),
    .B(_10997_),
    .ZN(_10998_));
 XNOR2_X1 _20672_ (.A(_10995_),
    .B(_10998_),
    .ZN(_10999_));
 MUX2_X1 _20673_ (.A(_10994_),
    .B(_10999_),
    .S(_10958_),
    .Z(_00661_));
 XOR2_X1 _20674_ (.A(_17076_),
    .B(_16972_),
    .Z(_11000_));
 XNOR2_X1 _20675_ (.A(_09603_),
    .B(_09685_),
    .ZN(_11001_));
 XNOR2_X1 _20676_ (.A(_11001_),
    .B(_09984_),
    .ZN(_11002_));
 XNOR2_X1 _20677_ (.A(_09372_),
    .B(_09258_),
    .ZN(_11003_));
 XNOR2_X1 _20678_ (.A(_11002_),
    .B(_11003_),
    .ZN(_11004_));
 XNOR2_X1 _20679_ (.A(_11004_),
    .B(_17076_),
    .ZN(_11005_));
 MUX2_X1 _20680_ (.A(_11000_),
    .B(_11005_),
    .S(_10958_),
    .Z(_00662_));
 XOR2_X1 _20681_ (.A(_17077_),
    .B(_16973_),
    .Z(_11006_));
 XNOR2_X1 _20682_ (.A(_09534_),
    .B(_10980_),
    .ZN(_11007_));
 XNOR2_X1 _20683_ (.A(_11007_),
    .B(_09836_),
    .ZN(_11008_));
 XOR2_X1 _20684_ (.A(_10954_),
    .B(_10060_),
    .Z(_11009_));
 XNOR2_X1 _20685_ (.A(_11008_),
    .B(_11009_),
    .ZN(_11010_));
 XNOR2_X1 _20686_ (.A(_11010_),
    .B(_10307_),
    .ZN(_11011_));
 INV_X1 _20687_ (.A(_17077_),
    .ZN(_11012_));
 XNOR2_X1 _20688_ (.A(_11011_),
    .B(_11012_),
    .ZN(_11013_));
 MUX2_X1 _20689_ (.A(_11006_),
    .B(_11013_),
    .S(_10958_),
    .Z(_00663_));
 XOR2_X1 _20690_ (.A(_17079_),
    .B(_16975_),
    .Z(_11014_));
 XNOR2_X1 _20691_ (.A(_09914_),
    .B(_10824_),
    .ZN(_11015_));
 XNOR2_X1 _20692_ (.A(_10960_),
    .B(_11015_),
    .ZN(_11016_));
 XOR2_X1 _20693_ (.A(_10181_),
    .B(_10119_),
    .Z(_11017_));
 XNOR2_X1 _20694_ (.A(_11017_),
    .B(_10542_),
    .ZN(_11018_));
 XNOR2_X1 _20695_ (.A(_11016_),
    .B(_11018_),
    .ZN(_11019_));
 XNOR2_X1 _20696_ (.A(_11019_),
    .B(_17079_),
    .ZN(_11020_));
 MUX2_X1 _20697_ (.A(_11014_),
    .B(_11020_),
    .S(_10958_),
    .Z(_00664_));
 XOR2_X1 _20698_ (.A(_16976_),
    .B(_17080_),
    .Z(_11021_));
 XNOR2_X1 _20699_ (.A(_10485_),
    .B(_10119_),
    .ZN(_11022_));
 XNOR2_X1 _20700_ (.A(_11022_),
    .B(_10770_),
    .ZN(_11023_));
 XNOR2_X1 _20701_ (.A(_10237_),
    .B(_01052_),
    .ZN(_11024_));
 XNOR2_X1 _20702_ (.A(_10371_),
    .B(_11024_),
    .ZN(_11025_));
 XNOR2_X1 _20703_ (.A(_11023_),
    .B(_11025_),
    .ZN(_11026_));
 BUF_X2 _20704_ (.A(_09039_),
    .Z(_11027_));
 MUX2_X1 _20705_ (.A(_11021_),
    .B(_11026_),
    .S(_11027_),
    .Z(_00665_));
 XOR2_X1 _20706_ (.A(_16977_),
    .B(_17081_),
    .Z(_11028_));
 XOR2_X1 _20707_ (.A(_10371_),
    .B(_10604_),
    .Z(_11029_));
 XNOR2_X1 _20708_ (.A(_11029_),
    .B(_10924_),
    .ZN(_11030_));
 XNOR2_X1 _20709_ (.A(_10431_),
    .B(_01053_),
    .ZN(_11031_));
 XNOR2_X1 _20710_ (.A(_11031_),
    .B(_10705_),
    .ZN(_11032_));
 XNOR2_X1 _20711_ (.A(_11030_),
    .B(_11032_),
    .ZN(_11033_));
 MUX2_X1 _20712_ (.A(_11028_),
    .B(_11033_),
    .S(_11027_),
    .Z(_00666_));
 XOR2_X1 _20713_ (.A(_17082_),
    .B(_16978_),
    .Z(_11034_));
 XNOR2_X1 _20714_ (.A(_10651_),
    .B(_10871_),
    .ZN(_11035_));
 XNOR2_X1 _20715_ (.A(_11035_),
    .B(_10979_),
    .ZN(_11036_));
 XNOR2_X1 _20716_ (.A(_11036_),
    .B(_09035_),
    .ZN(_11037_));
 XNOR2_X1 _20717_ (.A(_11037_),
    .B(_17082_),
    .ZN(_11038_));
 MUX2_X1 _20718_ (.A(_11034_),
    .B(_11038_),
    .S(_11027_),
    .Z(_00667_));
 CLKBUF_X2 _20719_ (.A(_17083_),
    .Z(_11039_));
 BUF_X2 _20720_ (.A(_11039_),
    .Z(_11040_));
 XOR2_X1 _20721_ (.A(_16979_),
    .B(_11040_),
    .Z(_11041_));
 XOR2_X1 _20722_ (.A(_10997_),
    .B(_01054_),
    .Z(_11042_));
 XNOR2_X1 _20723_ (.A(_06677_),
    .B(_08811_),
    .ZN(_11043_));
 XNOR2_X1 _20724_ (.A(_11043_),
    .B(_09147_),
    .ZN(_11044_));
 XNOR2_X1 _20725_ (.A(_11042_),
    .B(_11044_),
    .ZN(_11045_));
 MUX2_X1 _20726_ (.A(_11041_),
    .B(_11045_),
    .S(_11027_),
    .Z(_00628_));
 BUF_X2 _20727_ (.A(_17084_),
    .Z(_11046_));
 XOR2_X1 _20728_ (.A(_16980_),
    .B(_11046_),
    .Z(_11047_));
 XOR2_X1 _20729_ (.A(_09758_),
    .B(_01055_),
    .Z(_11048_));
 XNOR2_X1 _20730_ (.A(_11003_),
    .B(_11048_),
    .ZN(_11049_));
 XNOR2_X1 _20731_ (.A(_10997_),
    .B(_08814_),
    .ZN(_11050_));
 XNOR2_X1 _20732_ (.A(_11049_),
    .B(_11050_),
    .ZN(_11051_));
 MUX2_X1 _20733_ (.A(_11047_),
    .B(_11051_),
    .S(_11027_),
    .Z(_00629_));
 XOR2_X1 _20734_ (.A(_17085_),
    .B(_16981_),
    .Z(_11052_));
 XOR2_X1 _20735_ (.A(_09534_),
    .B(_09685_),
    .Z(_11053_));
 XNOR2_X1 _20736_ (.A(_11053_),
    .B(_09448_),
    .ZN(_11054_));
 XNOR2_X1 _20737_ (.A(_11054_),
    .B(_09984_),
    .ZN(_11055_));
 XNOR2_X1 _20738_ (.A(_11055_),
    .B(_17085_),
    .ZN(_11056_));
 MUX2_X1 _20739_ (.A(_11052_),
    .B(_11056_),
    .S(_11027_),
    .Z(_00630_));
 XOR2_X1 _20740_ (.A(_17086_),
    .B(_16982_),
    .Z(_11057_));
 XNOR2_X1 _20741_ (.A(_09987_),
    .B(_09914_),
    .ZN(_11058_));
 XNOR2_X1 _20742_ (.A(_11058_),
    .B(_10307_),
    .ZN(_11059_));
 XOR2_X1 _20743_ (.A(_11007_),
    .B(_10060_),
    .Z(_11060_));
 XNOR2_X1 _20744_ (.A(_11059_),
    .B(_11060_),
    .ZN(_11061_));
 INV_X1 _20745_ (.A(_17086_),
    .ZN(_11062_));
 XNOR2_X1 _20746_ (.A(_11061_),
    .B(_11062_),
    .ZN(_11063_));
 MUX2_X1 _20747_ (.A(_11057_),
    .B(_11063_),
    .S(_11027_),
    .Z(_00631_));
 XOR2_X1 _20748_ (.A(_17087_),
    .B(_16983_),
    .Z(_11064_));
 XNOR2_X1 _20749_ (.A(_10065_),
    .B(_11015_),
    .ZN(_11065_));
 XNOR2_X1 _20750_ (.A(_10119_),
    .B(_10237_),
    .ZN(_11066_));
 XNOR2_X1 _20751_ (.A(_11066_),
    .B(_10542_),
    .ZN(_11067_));
 XNOR2_X1 _20752_ (.A(_11065_),
    .B(_11067_),
    .ZN(_11068_));
 XNOR2_X1 _20753_ (.A(_11068_),
    .B(_17087_),
    .ZN(_11069_));
 MUX2_X1 _20754_ (.A(_11064_),
    .B(_11069_),
    .S(_11027_),
    .Z(_00632_));
 XOR2_X1 _20755_ (.A(_16984_),
    .B(_17088_),
    .Z(_11070_));
 XNOR2_X1 _20756_ (.A(_10431_),
    .B(_01056_),
    .ZN(_11071_));
 XNOR2_X1 _20757_ (.A(_11071_),
    .B(_10371_),
    .ZN(_11072_));
 XOR2_X1 _20758_ (.A(_10238_),
    .B(_10770_),
    .Z(_11073_));
 XNOR2_X1 _20759_ (.A(_11072_),
    .B(_11073_),
    .ZN(_11074_));
 MUX2_X1 _20760_ (.A(_11070_),
    .B(_11074_),
    .S(_11027_),
    .Z(_00633_));
 XOR2_X1 _20761_ (.A(_16986_),
    .B(_17090_),
    .Z(_11075_));
 XOR2_X1 _20762_ (.A(_10651_),
    .B(_10705_),
    .Z(_11076_));
 XNOR2_X1 _20763_ (.A(_10924_),
    .B(_01057_),
    .ZN(_11077_));
 XNOR2_X1 _20764_ (.A(_11076_),
    .B(_11077_),
    .ZN(_11078_));
 XNOR2_X1 _20765_ (.A(_11078_),
    .B(_10486_),
    .ZN(_11079_));
 MUX2_X1 _20766_ (.A(_11075_),
    .B(_11079_),
    .S(_11027_),
    .Z(_00634_));
 XOR2_X1 _20767_ (.A(_17091_),
    .B(_16987_),
    .Z(_11080_));
 XNOR2_X1 _20768_ (.A(_10652_),
    .B(_10872_),
    .ZN(_11081_));
 XNOR2_X1 _20769_ (.A(_11081_),
    .B(_09035_),
    .ZN(_11082_));
 XNOR2_X1 _20770_ (.A(_11082_),
    .B(_17091_),
    .ZN(_11083_));
 BUF_X2 _20771_ (.A(_09039_),
    .Z(_11084_));
 MUX2_X1 _20772_ (.A(_11080_),
    .B(_11083_),
    .S(_11084_),
    .Z(_00635_));
 XOR2_X1 _20773_ (.A(_17163_),
    .B(_16988_),
    .Z(_11085_));
 INV_X1 _20774_ (.A(_16739_),
    .ZN(_11086_));
 AND2_X1 _20775_ (.A1(_11086_),
    .A2(_16740_),
    .ZN(_11087_));
 CLKBUF_X2 _20776_ (.A(_11087_),
    .Z(_11088_));
 INV_X1 _20777_ (.A(_16741_),
    .ZN(_11089_));
 NOR2_X1 _20778_ (.A1(_11089_),
    .A2(_16742_),
    .ZN(_11090_));
 CLKBUF_X2 _20779_ (.A(_11090_),
    .Z(_11091_));
 AND2_X1 _20780_ (.A1(_11088_),
    .A2(_11091_),
    .ZN(_11092_));
 BUF_X2 _20781_ (.A(_11092_),
    .Z(_11093_));
 NOR2_X1 _20782_ (.A1(_16737_),
    .A2(_16738_),
    .ZN(_11094_));
 CLKBUF_X2 _20783_ (.A(_16735_),
    .Z(_11095_));
 AND2_X1 _20784_ (.A1(_11094_),
    .A2(_11095_),
    .ZN(_11096_));
 INV_X1 _20785_ (.A(_16737_),
    .ZN(_11097_));
 NOR2_X2 _20786_ (.A1(_11097_),
    .A2(_16738_),
    .ZN(_11098_));
 CLKBUF_X2 _20787_ (.A(_11098_),
    .Z(_11099_));
 BUF_X2 _20788_ (.A(_11099_),
    .Z(_11100_));
 OAI21_X1 _20789_ (.A(_11093_),
    .B1(_11096_),
    .B2(_11100_),
    .ZN(_11101_));
 AND2_X1 _20790_ (.A1(_16740_),
    .A2(_16739_),
    .ZN(_11102_));
 AND2_X1 _20791_ (.A1(_11090_),
    .A2(_11102_),
    .ZN(_11103_));
 AND2_X1 _20792_ (.A1(_16736_),
    .A2(_16735_),
    .ZN(_11104_));
 AND2_X2 _20793_ (.A1(_11104_),
    .A2(_11094_),
    .ZN(_11105_));
 NAND2_X1 _20794_ (.A1(_11103_),
    .A2(_11105_),
    .ZN(_11106_));
 INV_X1 _20795_ (.A(_11103_),
    .ZN(_11107_));
 INV_X1 _20796_ (.A(_16736_),
    .ZN(_11108_));
 CLKBUF_X2 _20797_ (.A(_11108_),
    .Z(_11109_));
 AND2_X1 _20798_ (.A1(_11094_),
    .A2(_11109_),
    .ZN(_11110_));
 INV_X1 _20799_ (.A(_11110_),
    .ZN(_11111_));
 OAI21_X1 _20800_ (.A(_11106_),
    .B1(_11107_),
    .B2(_11111_),
    .ZN(_11112_));
 INV_X1 _20801_ (.A(_16738_),
    .ZN(_11113_));
 NOR2_X2 _20802_ (.A1(_11113_),
    .A2(_16737_),
    .ZN(_11114_));
 CLKBUF_X2 _20803_ (.A(_11104_),
    .Z(_11115_));
 AND2_X2 _20804_ (.A1(_11114_),
    .A2(_11115_),
    .ZN(_11116_));
 INV_X1 _20805_ (.A(_11116_),
    .ZN(_11117_));
 NOR2_X2 _20806_ (.A1(_11108_),
    .A2(_16735_),
    .ZN(_11118_));
 AND2_X1 _20807_ (.A1(_16737_),
    .A2(_16738_),
    .ZN(_11119_));
 AND2_X1 _20808_ (.A1(_11118_),
    .A2(_11119_),
    .ZN(_11120_));
 BUF_X2 _20809_ (.A(_11120_),
    .Z(_11121_));
 INV_X1 _20810_ (.A(_11121_),
    .ZN(_11122_));
 AOI21_X1 _20811_ (.A(_11107_),
    .B1(_11117_),
    .B2(_11122_),
    .ZN(_11123_));
 INV_X1 _20812_ (.A(_16735_),
    .ZN(_11124_));
 NOR2_X2 _20813_ (.A1(_11124_),
    .A2(_16736_),
    .ZN(_11125_));
 CLKBUF_X2 _20814_ (.A(_11119_),
    .Z(_11126_));
 AND2_X1 _20815_ (.A1(_11125_),
    .A2(_11126_),
    .ZN(_11127_));
 BUF_X2 _20816_ (.A(_11127_),
    .Z(_11128_));
 BUF_X2 _20817_ (.A(_11103_),
    .Z(_11129_));
 AND2_X1 _20818_ (.A1(_11128_),
    .A2(_11129_),
    .ZN(_11130_));
 OR2_X1 _20819_ (.A1(_11123_),
    .A2(_11130_),
    .ZN(_11131_));
 NOR2_X1 _20820_ (.A1(_11124_),
    .A2(_16738_),
    .ZN(_11132_));
 AND2_X1 _20821_ (.A1(_11132_),
    .A2(_16737_),
    .ZN(_11133_));
 AOI211_X1 _20822_ (.A(_11112_),
    .B(_11131_),
    .C1(_11129_),
    .C2(_11133_),
    .ZN(_11134_));
 NOR2_X2 _20823_ (.A1(_16740_),
    .A2(_16739_),
    .ZN(_11135_));
 AND2_X1 _20824_ (.A1(_11091_),
    .A2(_11135_),
    .ZN(_11136_));
 BUF_X2 _20825_ (.A(_11136_),
    .Z(_11137_));
 AND2_X1 _20826_ (.A1(_11126_),
    .A2(_11109_),
    .ZN(_11138_));
 CLKBUF_X2 _20827_ (.A(_11138_),
    .Z(_11139_));
 OAI21_X1 _20828_ (.A(_11137_),
    .B1(_11121_),
    .B2(_11139_),
    .ZN(_11140_));
 CLKBUF_X2 _20829_ (.A(_11114_),
    .Z(_11141_));
 BUF_X2 _20830_ (.A(_11095_),
    .Z(_11142_));
 BUF_X2 _20831_ (.A(_11135_),
    .Z(_11143_));
 NAND4_X1 _20832_ (.A1(_11141_),
    .A2(_11091_),
    .A3(_11142_),
    .A4(_11143_),
    .ZN(_11144_));
 NAND2_X1 _20833_ (.A1(_11140_),
    .A2(_11144_),
    .ZN(_11145_));
 INV_X1 _20834_ (.A(_11145_),
    .ZN(_11146_));
 NOR2_X1 _20835_ (.A1(_11086_),
    .A2(_16740_),
    .ZN(_11147_));
 AND2_X2 _20836_ (.A1(_11090_),
    .A2(_11147_),
    .ZN(_11148_));
 BUF_X2 _20837_ (.A(_11148_),
    .Z(_11149_));
 CLKBUF_X2 _20838_ (.A(_16736_),
    .Z(_11150_));
 AND2_X1 _20839_ (.A1(_11098_),
    .A2(_11150_),
    .ZN(_11151_));
 BUF_X2 _20840_ (.A(_11151_),
    .Z(_11152_));
 BUF_X2 _20841_ (.A(_11094_),
    .Z(_11153_));
 INV_X1 _20842_ (.A(_11153_),
    .ZN(_11154_));
 CLKBUF_X2 _20843_ (.A(_11118_),
    .Z(_11155_));
 NOR2_X1 _20844_ (.A1(_11154_),
    .A2(_11155_),
    .ZN(_11156_));
 OAI21_X1 _20845_ (.A(_11149_),
    .B1(_11152_),
    .B2(_11156_),
    .ZN(_11157_));
 NOR2_X2 _20846_ (.A1(_16736_),
    .A2(_16735_),
    .ZN(_11158_));
 AND2_X1 _20847_ (.A1(_11098_),
    .A2(_11158_),
    .ZN(_11159_));
 CLKBUF_X2 _20848_ (.A(_11110_),
    .Z(_11160_));
 OAI21_X1 _20849_ (.A(_11137_),
    .B1(_11159_),
    .B2(_11160_),
    .ZN(_11161_));
 AND2_X1 _20850_ (.A1(_11114_),
    .A2(_11095_),
    .ZN(_11162_));
 AND2_X1 _20851_ (.A1(_11115_),
    .A2(_11126_),
    .ZN(_11163_));
 OAI21_X1 _20852_ (.A(_11149_),
    .B1(_11162_),
    .B2(_11163_),
    .ZN(_11164_));
 AND4_X1 _20853_ (.A1(_11146_),
    .A2(_11157_),
    .A3(_11161_),
    .A4(_11164_),
    .ZN(_11165_));
 NOR3_X1 _20854_ (.A1(_11118_),
    .A2(_16737_),
    .A3(_11113_),
    .ZN(_11166_));
 OAI21_X1 _20855_ (.A(_11093_),
    .B1(_11166_),
    .B2(_11121_),
    .ZN(_11167_));
 AND4_X1 _20856_ (.A1(_11101_),
    .A2(_11134_),
    .A3(_11165_),
    .A4(_11167_),
    .ZN(_11168_));
 INV_X1 _20857_ (.A(_11114_),
    .ZN(_11169_));
 NOR2_X2 _20858_ (.A1(_16742_),
    .A2(_16741_),
    .ZN(_11170_));
 AND2_X1 _20859_ (.A1(_11170_),
    .A2(_11135_),
    .ZN(_11171_));
 INV_X1 _20860_ (.A(_11171_),
    .ZN(_11172_));
 CLKBUF_X2 _20861_ (.A(_11124_),
    .Z(_11173_));
 AOI211_X1 _20862_ (.A(_11169_),
    .B(_11172_),
    .C1(_11109_),
    .C2(_11173_),
    .ZN(_11174_));
 CLKBUF_X2 _20863_ (.A(_11171_),
    .Z(_11175_));
 NAND2_X1 _20864_ (.A1(_11152_),
    .A2(_11175_),
    .ZN(_11176_));
 AND2_X2 _20865_ (.A1(_11125_),
    .A2(_11098_),
    .ZN(_11177_));
 INV_X1 _20866_ (.A(_11177_),
    .ZN(_11178_));
 OAI21_X1 _20867_ (.A(_11176_),
    .B1(_11178_),
    .B2(_11172_),
    .ZN(_11179_));
 AND2_X1 _20868_ (.A1(_11094_),
    .A2(_11150_),
    .ZN(_11180_));
 BUF_X2 _20869_ (.A(_11180_),
    .Z(_11181_));
 AND2_X1 _20870_ (.A1(_11175_),
    .A2(_11181_),
    .ZN(_11182_));
 INV_X1 _20871_ (.A(_11104_),
    .ZN(_11183_));
 CLKBUF_X2 _20872_ (.A(_11183_),
    .Z(_11184_));
 CLKBUF_X2 _20873_ (.A(_11126_),
    .Z(_11185_));
 INV_X2 _20874_ (.A(_11158_),
    .ZN(_11186_));
 AND4_X1 _20875_ (.A1(_11184_),
    .A2(_11175_),
    .A3(_11185_),
    .A4(_11186_),
    .ZN(_11187_));
 NOR4_X1 _20876_ (.A1(_11174_),
    .A2(_11179_),
    .A3(_11182_),
    .A4(_11187_),
    .ZN(_11188_));
 BUF_X2 _20877_ (.A(_11158_),
    .Z(_11189_));
 NOR2_X2 _20878_ (.A1(_11154_),
    .A2(_11189_),
    .ZN(_11190_));
 AND2_X1 _20879_ (.A1(_11102_),
    .A2(_11170_),
    .ZN(_11191_));
 AND2_X1 _20880_ (.A1(_11190_),
    .A2(_11191_),
    .ZN(_11192_));
 CLKBUF_X2 _20881_ (.A(_11170_),
    .Z(_11193_));
 BUF_X2 _20882_ (.A(_11099_),
    .Z(_11194_));
 CLKBUF_X2 _20883_ (.A(_11102_),
    .Z(_11195_));
 AND4_X1 _20884_ (.A1(_11193_),
    .A2(_11194_),
    .A3(_11155_),
    .A4(_11195_),
    .ZN(_11196_));
 OR2_X1 _20885_ (.A1(_11192_),
    .A2(_11196_),
    .ZN(_11197_));
 AND2_X1 _20886_ (.A1(_11163_),
    .A2(_11191_),
    .ZN(_11198_));
 CLKBUF_X2 _20887_ (.A(_11191_),
    .Z(_11199_));
 AND3_X1 _20888_ (.A1(_11199_),
    .A2(_11189_),
    .A3(_11141_),
    .ZN(_11200_));
 AND2_X1 _20889_ (.A1(_11139_),
    .A2(_11199_),
    .ZN(_11201_));
 NOR4_X1 _20890_ (.A1(_11197_),
    .A2(_11198_),
    .A3(_11200_),
    .A4(_11201_),
    .ZN(_11202_));
 INV_X1 _20891_ (.A(_11125_),
    .ZN(_11203_));
 AND2_X1 _20892_ (.A1(_11166_),
    .A2(_11203_),
    .ZN(_11204_));
 AND2_X1 _20893_ (.A1(_11147_),
    .A2(_11170_),
    .ZN(_11205_));
 AND2_X1 _20894_ (.A1(_11204_),
    .A2(_11205_),
    .ZN(_11206_));
 BUF_X2 _20895_ (.A(_11205_),
    .Z(_11207_));
 NAND4_X1 _20896_ (.A1(_11207_),
    .A2(_11184_),
    .A3(_11186_),
    .A4(_11100_),
    .ZN(_11208_));
 INV_X1 _20897_ (.A(_11205_),
    .ZN(_11209_));
 INV_X1 _20898_ (.A(_11181_),
    .ZN(_11210_));
 OAI21_X1 _20899_ (.A(_11208_),
    .B1(_11209_),
    .B2(_11210_),
    .ZN(_11211_));
 NOR2_X1 _20900_ (.A1(_11206_),
    .A2(_11211_),
    .ZN(_11212_));
 AND2_X1 _20901_ (.A1(_11088_),
    .A2(_11170_),
    .ZN(_11213_));
 INV_X1 _20902_ (.A(_11213_),
    .ZN(_11214_));
 AND2_X2 _20903_ (.A1(_11126_),
    .A2(_11158_),
    .ZN(_11215_));
 INV_X1 _20904_ (.A(_11215_),
    .ZN(_11216_));
 AND2_X1 _20905_ (.A1(_11126_),
    .A2(_11150_),
    .ZN(_11217_));
 INV_X1 _20906_ (.A(_11217_),
    .ZN(_11218_));
 AOI21_X1 _20907_ (.A(_11214_),
    .B1(_11216_),
    .B2(_11218_),
    .ZN(_11219_));
 AND2_X1 _20908_ (.A1(_11183_),
    .A2(_11099_),
    .ZN(_11220_));
 CLKBUF_X2 _20909_ (.A(_11213_),
    .Z(_11221_));
 AND3_X1 _20910_ (.A1(_11220_),
    .A2(_11186_),
    .A3(_11221_),
    .ZN(_11222_));
 NOR2_X1 _20911_ (.A1(_11154_),
    .A2(_11115_),
    .ZN(_11223_));
 AND2_X1 _20912_ (.A1(_11221_),
    .A2(_11223_),
    .ZN(_11224_));
 AND2_X1 _20913_ (.A1(_11186_),
    .A2(_11114_),
    .ZN(_11225_));
 AND2_X1 _20914_ (.A1(_11221_),
    .A2(_11225_),
    .ZN(_11226_));
 NOR4_X1 _20915_ (.A1(_11219_),
    .A2(_11222_),
    .A3(_11224_),
    .A4(_11226_),
    .ZN(_11227_));
 AND4_X1 _20916_ (.A1(_11188_),
    .A2(_11202_),
    .A3(_11212_),
    .A4(_11227_),
    .ZN(_11228_));
 INV_X1 _20917_ (.A(_11098_),
    .ZN(_11229_));
 NOR2_X1 _20918_ (.A1(_11229_),
    .A2(_11118_),
    .ZN(_11230_));
 AND2_X1 _20919_ (.A1(_11089_),
    .A2(_16742_),
    .ZN(_11231_));
 AND2_X1 _20920_ (.A1(_11231_),
    .A2(_11135_),
    .ZN(_11232_));
 NAND2_X1 _20921_ (.A1(_11230_),
    .A2(_11232_),
    .ZN(_11233_));
 BUF_X2 _20922_ (.A(_11232_),
    .Z(_11234_));
 BUF_X2 _20923_ (.A(_11217_),
    .Z(_11235_));
 OAI21_X1 _20924_ (.A(_11234_),
    .B1(_11128_),
    .B2(_11235_),
    .ZN(_11236_));
 CLKBUF_X2 _20925_ (.A(_11231_),
    .Z(_11237_));
 CLKBUF_X2 _20926_ (.A(_11237_),
    .Z(_11238_));
 BUF_X2 _20927_ (.A(_11153_),
    .Z(_11239_));
 NAND4_X1 _20928_ (.A1(_11238_),
    .A2(_11173_),
    .A3(_11143_),
    .A4(_11239_),
    .ZN(_11240_));
 NAND4_X1 _20929_ (.A1(_11238_),
    .A2(_11141_),
    .A3(_11142_),
    .A4(_11143_),
    .ZN(_11241_));
 AND4_X1 _20930_ (.A1(_11233_),
    .A2(_11236_),
    .A3(_11240_),
    .A4(_11241_),
    .ZN(_11242_));
 AND2_X1 _20931_ (.A1(_11231_),
    .A2(_11102_),
    .ZN(_11243_));
 AND2_X1 _20932_ (.A1(_11230_),
    .A2(_11243_),
    .ZN(_11244_));
 INV_X1 _20933_ (.A(_11244_),
    .ZN(_11245_));
 NAND3_X1 _20934_ (.A1(_11215_),
    .A2(_11238_),
    .A3(_11195_),
    .ZN(_11246_));
 BUF_X2 _20935_ (.A(_11243_),
    .Z(_11247_));
 AND2_X2 _20936_ (.A1(_11158_),
    .A2(_11094_),
    .ZN(_11248_));
 OAI21_X1 _20937_ (.A(_11247_),
    .B1(_11248_),
    .B2(_11181_),
    .ZN(_11249_));
 AND3_X1 _20938_ (.A1(_11245_),
    .A2(_11246_),
    .A3(_11249_),
    .ZN(_11250_));
 AND2_X1 _20939_ (.A1(_11231_),
    .A2(_11147_),
    .ZN(_11251_));
 BUF_X2 _20940_ (.A(_11251_),
    .Z(_11252_));
 AND3_X1 _20941_ (.A1(_11252_),
    .A2(_11186_),
    .A3(_11223_),
    .ZN(_11253_));
 AOI21_X1 _20942_ (.A(_11253_),
    .B1(_11235_),
    .B2(_11252_),
    .ZN(_11254_));
 BUF_X2 _20943_ (.A(_11088_),
    .Z(_11255_));
 OAI211_X1 _20944_ (.A(_11255_),
    .B(_11238_),
    .C1(_11163_),
    .C2(_11139_),
    .ZN(_11256_));
 NAND4_X1 _20945_ (.A1(_11255_),
    .A2(_11238_),
    .A3(_11125_),
    .A4(_11141_),
    .ZN(_11257_));
 AND2_X1 _20946_ (.A1(_11087_),
    .A2(_11231_),
    .ZN(_11258_));
 BUF_X2 _20947_ (.A(_11258_),
    .Z(_11259_));
 NAND2_X1 _20948_ (.A1(_11259_),
    .A2(_11159_),
    .ZN(_11260_));
 AND3_X1 _20949_ (.A1(_11256_),
    .A2(_11257_),
    .A3(_11260_),
    .ZN(_11261_));
 AND4_X1 _20950_ (.A1(_11242_),
    .A2(_11250_),
    .A3(_11254_),
    .A4(_11261_),
    .ZN(_11262_));
 AND2_X1 _20951_ (.A1(_16742_),
    .A2(_16741_),
    .ZN(_11263_));
 AND2_X2 _20952_ (.A1(_11147_),
    .A2(_11263_),
    .ZN(_11264_));
 BUF_X2 _20953_ (.A(_11264_),
    .Z(_11265_));
 INV_X1 _20954_ (.A(_11128_),
    .ZN(_11266_));
 AND2_X1 _20955_ (.A1(_11118_),
    .A2(_11153_),
    .ZN(_11267_));
 INV_X1 _20956_ (.A(_11267_),
    .ZN(_11268_));
 NAND3_X1 _20957_ (.A1(_11178_),
    .A2(_11266_),
    .A3(_11268_),
    .ZN(_11269_));
 INV_X1 _20958_ (.A(_11118_),
    .ZN(_11270_));
 AOI21_X1 _20959_ (.A(_11113_),
    .B1(_11270_),
    .B2(_16737_),
    .ZN(_11271_));
 OAI21_X1 _20960_ (.A(_11265_),
    .B1(_11269_),
    .B2(_11271_),
    .ZN(_11272_));
 NOR2_X1 _20961_ (.A1(_11169_),
    .A2(_11125_),
    .ZN(_11273_));
 AND2_X2 _20962_ (.A1(_11088_),
    .A2(_11263_),
    .ZN(_11274_));
 AND2_X1 _20963_ (.A1(_11273_),
    .A2(_11274_),
    .ZN(_11275_));
 INV_X1 _20964_ (.A(_11274_),
    .ZN(_11276_));
 INV_X1 _20965_ (.A(_11105_),
    .ZN(_11277_));
 INV_X1 _20966_ (.A(_11248_),
    .ZN(_11278_));
 NAND2_X1 _20967_ (.A1(_11277_),
    .A2(_11278_),
    .ZN(_11279_));
 INV_X1 _20968_ (.A(_11279_),
    .ZN(_11280_));
 AND2_X1 _20969_ (.A1(_11098_),
    .A2(_11109_),
    .ZN(_11281_));
 BUF_X2 _20970_ (.A(_11281_),
    .Z(_11282_));
 INV_X1 _20971_ (.A(_11282_),
    .ZN(_11283_));
 AOI21_X1 _20972_ (.A(_11276_),
    .B1(_11280_),
    .B2(_11283_),
    .ZN(_11284_));
 BUF_X2 _20973_ (.A(_11274_),
    .Z(_11285_));
 AND2_X1 _20974_ (.A1(_11126_),
    .A2(_11095_),
    .ZN(_11286_));
 AOI211_X1 _20975_ (.A(_11275_),
    .B(_11284_),
    .C1(_11285_),
    .C2(_11286_),
    .ZN(_11287_));
 CLKBUF_X2 _20976_ (.A(_11263_),
    .Z(_11288_));
 AND4_X1 _20977_ (.A1(_11143_),
    .A2(_11155_),
    .A3(_11239_),
    .A4(_11288_),
    .ZN(_11289_));
 AND2_X1 _20978_ (.A1(_11263_),
    .A2(_11135_),
    .ZN(_11290_));
 CLKBUF_X2 _20979_ (.A(_11290_),
    .Z(_11291_));
 INV_X1 _20980_ (.A(_11291_),
    .ZN(_11292_));
 INV_X1 _20981_ (.A(_11138_),
    .ZN(_11293_));
 AOI21_X1 _20982_ (.A(_11292_),
    .B1(_11122_),
    .B2(_11293_),
    .ZN(_11294_));
 BUF_X2 _20983_ (.A(_11291_),
    .Z(_11295_));
 AOI211_X1 _20984_ (.A(_11289_),
    .B(_11294_),
    .C1(_11162_),
    .C2(_11295_),
    .ZN(_11296_));
 AND2_X2 _20985_ (.A1(_11102_),
    .A2(_11263_),
    .ZN(_11297_));
 NAND2_X1 _20986_ (.A1(_11159_),
    .A2(_11297_),
    .ZN(_11298_));
 BUF_X2 _20987_ (.A(_11297_),
    .Z(_11299_));
 NOR2_X1 _20988_ (.A1(_11113_),
    .A2(_16736_),
    .ZN(_11300_));
 AND2_X2 _20989_ (.A1(_11300_),
    .A2(_11097_),
    .ZN(_11301_));
 BUF_X2 _20990_ (.A(_11301_),
    .Z(_11302_));
 AND2_X1 _20991_ (.A1(_11114_),
    .A2(_11150_),
    .ZN(_11303_));
 BUF_X2 _20992_ (.A(_11303_),
    .Z(_11304_));
 OAI21_X1 _20993_ (.A(_11299_),
    .B1(_11302_),
    .B2(_11304_),
    .ZN(_11305_));
 OAI211_X1 _20994_ (.A(_11299_),
    .B(_11239_),
    .C1(_11150_),
    .C2(_11142_),
    .ZN(_11306_));
 NAND3_X1 _20995_ (.A1(_11297_),
    .A2(_11185_),
    .A3(_11155_),
    .ZN(_11307_));
 AND4_X1 _20996_ (.A1(_11298_),
    .A2(_11305_),
    .A3(_11306_),
    .A4(_11307_),
    .ZN(_11308_));
 AND4_X1 _20997_ (.A1(_11272_),
    .A2(_11287_),
    .A3(_11296_),
    .A4(_11308_),
    .ZN(_11309_));
 NAND4_X1 _20998_ (.A1(_11168_),
    .A2(_11228_),
    .A3(_11262_),
    .A4(_11309_),
    .ZN(_11310_));
 AND2_X2 _20999_ (.A1(_11171_),
    .A2(_11248_),
    .ZN(_11311_));
 NOR2_X2 _21000_ (.A1(_11310_),
    .A2(_11311_),
    .ZN(_11312_));
 INV_X1 _21001_ (.A(_16749_),
    .ZN(_11313_));
 NOR2_X2 _21002_ (.A1(_11313_),
    .A2(_16750_),
    .ZN(_11314_));
 INV_X1 _21003_ (.A(_16747_),
    .ZN(_11315_));
 NOR2_X2 _21004_ (.A1(_11315_),
    .A2(_16748_),
    .ZN(_11316_));
 AND2_X1 _21005_ (.A1(_11314_),
    .A2(_11316_),
    .ZN(_11317_));
 CLKBUF_X2 _21006_ (.A(_11317_),
    .Z(_11318_));
 AND2_X2 _21007_ (.A1(_16744_),
    .A2(_16743_),
    .ZN(_11319_));
 NOR2_X2 _21008_ (.A1(_16745_),
    .A2(_16746_),
    .ZN(_11320_));
 AND2_X2 _21009_ (.A1(_11319_),
    .A2(_11320_),
    .ZN(_11321_));
 AND2_X1 _21010_ (.A1(_11318_),
    .A2(_11321_),
    .ZN(_11322_));
 INV_X1 _21011_ (.A(_11322_),
    .ZN(_11323_));
 INV_X1 _21012_ (.A(_11317_),
    .ZN(_11324_));
 INV_X1 _21013_ (.A(_16744_),
    .ZN(_11325_));
 AND2_X1 _21014_ (.A1(_11320_),
    .A2(_11325_),
    .ZN(_11326_));
 BUF_X2 _21015_ (.A(_11326_),
    .Z(_11327_));
 INV_X1 _21016_ (.A(_11327_),
    .ZN(_11328_));
 AND2_X1 _21017_ (.A1(_11315_),
    .A2(_16748_),
    .ZN(_11329_));
 AND2_X1 _21018_ (.A1(_11329_),
    .A2(_11314_),
    .ZN(_11330_));
 CLKBUF_X2 _21019_ (.A(_11330_),
    .Z(_11331_));
 INV_X1 _21020_ (.A(_16746_),
    .ZN(_11332_));
 NOR2_X2 _21021_ (.A1(_11332_),
    .A2(_16745_),
    .ZN(_11333_));
 CLKBUF_X2 _21022_ (.A(_11333_),
    .Z(_11334_));
 BUF_X2 _21023_ (.A(_16743_),
    .Z(_11335_));
 AND2_X1 _21024_ (.A1(_11334_),
    .A2(_11335_),
    .ZN(_11336_));
 NAND2_X1 _21025_ (.A1(_11331_),
    .A2(_11336_),
    .ZN(_11337_));
 BUF_X2 _21026_ (.A(_16744_),
    .Z(_11338_));
 OAI221_X1 _21027_ (.A(_11323_),
    .B1(_11324_),
    .B2(_11328_),
    .C1(_11337_),
    .C2(_11338_),
    .ZN(_11339_));
 AND2_X1 _21028_ (.A1(_11333_),
    .A2(_11319_),
    .ZN(_11340_));
 INV_X1 _21029_ (.A(_11340_),
    .ZN(_11341_));
 NOR2_X1 _21030_ (.A1(_16744_),
    .A2(_16743_),
    .ZN(_11342_));
 CLKBUF_X2 _21031_ (.A(_11342_),
    .Z(_11343_));
 AND2_X2 _21032_ (.A1(_11333_),
    .A2(_11343_),
    .ZN(_11344_));
 INV_X1 _21033_ (.A(_11344_),
    .ZN(_11345_));
 NAND2_X1 _21034_ (.A1(_11341_),
    .A2(_11345_),
    .ZN(_11346_));
 CLKBUF_X2 _21035_ (.A(_11331_),
    .Z(_11347_));
 AND2_X1 _21036_ (.A1(_11346_),
    .A2(_11347_),
    .ZN(_11348_));
 AND2_X1 _21037_ (.A1(_11313_),
    .A2(_16750_),
    .ZN(_11349_));
 NOR2_X1 _21038_ (.A1(_16748_),
    .A2(_16747_),
    .ZN(_11350_));
 CLKBUF_X2 _21039_ (.A(_11350_),
    .Z(_11351_));
 AND2_X1 _21040_ (.A1(_11349_),
    .A2(_11351_),
    .ZN(_11352_));
 CLKBUF_X2 _21041_ (.A(_11352_),
    .Z(_11353_));
 AND2_X1 _21042_ (.A1(_16745_),
    .A2(_16746_),
    .ZN(_11354_));
 INV_X1 _21043_ (.A(_11354_),
    .ZN(_11355_));
 NOR2_X1 _21044_ (.A1(_11355_),
    .A2(_11343_),
    .ZN(_11356_));
 AND2_X1 _21045_ (.A1(_11353_),
    .A2(_11356_),
    .ZN(_11357_));
 OR3_X1 _21046_ (.A1(_11339_),
    .A2(_11348_),
    .A3(_11357_),
    .ZN(_11358_));
 INV_X1 _21047_ (.A(_11333_),
    .ZN(_11359_));
 INV_X1 _21048_ (.A(_16743_),
    .ZN(_11360_));
 NOR2_X1 _21049_ (.A1(_11360_),
    .A2(_16744_),
    .ZN(_11361_));
 CLKBUF_X2 _21050_ (.A(_11361_),
    .Z(_11362_));
 NOR2_X1 _21051_ (.A1(_11359_),
    .A2(_11362_),
    .ZN(_11363_));
 CLKBUF_X2 _21052_ (.A(_11329_),
    .Z(_11364_));
 AND2_X1 _21053_ (.A1(_16750_),
    .A2(_16749_),
    .ZN(_11365_));
 AND2_X1 _21054_ (.A1(_11364_),
    .A2(_11365_),
    .ZN(_11366_));
 AND2_X1 _21055_ (.A1(_11363_),
    .A2(_11366_),
    .ZN(_11367_));
 BUF_X2 _21056_ (.A(_11349_),
    .Z(_11368_));
 AND2_X1 _21057_ (.A1(_11319_),
    .A2(_11354_),
    .ZN(_11369_));
 BUF_X2 _21058_ (.A(_11369_),
    .Z(_11370_));
 AND2_X2 _21059_ (.A1(_11354_),
    .A2(_11325_),
    .ZN(_11371_));
 OAI211_X1 _21060_ (.A(_11364_),
    .B(_11368_),
    .C1(_11370_),
    .C2(_11371_),
    .ZN(_11372_));
 BUF_X2 _21061_ (.A(_11334_),
    .Z(_11373_));
 NAND4_X1 _21062_ (.A1(_11364_),
    .A2(_11368_),
    .A3(_11362_),
    .A4(_11373_),
    .ZN(_11374_));
 NAND2_X1 _21063_ (.A1(_11372_),
    .A2(_11374_),
    .ZN(_11375_));
 INV_X1 _21064_ (.A(_16745_),
    .ZN(_11376_));
 NOR2_X1 _21065_ (.A1(_11376_),
    .A2(_16746_),
    .ZN(_11377_));
 INV_X1 _21066_ (.A(_11377_),
    .ZN(_11378_));
 NOR2_X1 _21067_ (.A1(_11325_),
    .A2(_16743_),
    .ZN(_11379_));
 NOR2_X2 _21068_ (.A1(_11378_),
    .A2(_11379_),
    .ZN(_11380_));
 AND2_X1 _21069_ (.A1(_16748_),
    .A2(_16747_),
    .ZN(_11381_));
 AND2_X2 _21070_ (.A1(_11349_),
    .A2(_11381_),
    .ZN(_11382_));
 AND2_X1 _21071_ (.A1(_11380_),
    .A2(_11382_),
    .ZN(_11383_));
 NOR4_X1 _21072_ (.A1(_11358_),
    .A2(_11367_),
    .A3(_11375_),
    .A4(_11383_),
    .ZN(_11384_));
 NOR2_X2 _21073_ (.A1(_16750_),
    .A2(_16749_),
    .ZN(_11385_));
 AND2_X2 _21074_ (.A1(_11381_),
    .A2(_11385_),
    .ZN(_11386_));
 INV_X1 _21075_ (.A(_11386_),
    .ZN(_11387_));
 INV_X1 _21076_ (.A(_11342_),
    .ZN(_11388_));
 CLKBUF_X2 _21077_ (.A(_11320_),
    .Z(_11389_));
 NAND2_X1 _21078_ (.A1(_11388_),
    .A2(_11389_),
    .ZN(_11390_));
 NOR2_X1 _21079_ (.A1(_11387_),
    .A2(_11390_),
    .ZN(_11391_));
 INV_X1 _21080_ (.A(_11391_),
    .ZN(_11392_));
 AND2_X1 _21081_ (.A1(_11389_),
    .A2(_11360_),
    .ZN(_11393_));
 OAI21_X1 _21082_ (.A(_11353_),
    .B1(_11336_),
    .B2(_11393_),
    .ZN(_11394_));
 CLKBUF_X2 _21083_ (.A(_11377_),
    .Z(_11395_));
 CLKBUF_X2 _21084_ (.A(_11395_),
    .Z(_11396_));
 NAND4_X1 _21085_ (.A1(_11368_),
    .A2(_11396_),
    .A3(_11319_),
    .A4(_11351_),
    .ZN(_11397_));
 AND2_X2 _21086_ (.A1(_11395_),
    .A2(_11343_),
    .ZN(_11398_));
 NAND2_X1 _21087_ (.A1(_11352_),
    .A2(_11398_),
    .ZN(_11399_));
 AND2_X2 _21088_ (.A1(_11395_),
    .A2(_11361_),
    .ZN(_11400_));
 NAND3_X1 _21089_ (.A1(_11400_),
    .A2(_11351_),
    .A3(_11368_),
    .ZN(_11401_));
 AND4_X1 _21090_ (.A1(_11394_),
    .A2(_11397_),
    .A3(_11399_),
    .A4(_11401_),
    .ZN(_11402_));
 BUF_X2 _21091_ (.A(_11318_),
    .Z(_11403_));
 OAI21_X1 _21092_ (.A(_11403_),
    .B1(_11336_),
    .B2(_11370_),
    .ZN(_11404_));
 AND2_X1 _21093_ (.A1(_11314_),
    .A2(_11381_),
    .ZN(_11405_));
 BUF_X2 _21094_ (.A(_11405_),
    .Z(_11406_));
 INV_X1 _21095_ (.A(_11319_),
    .ZN(_11407_));
 CLKBUF_X2 _21096_ (.A(_11407_),
    .Z(_11408_));
 AND2_X1 _21097_ (.A1(_11356_),
    .A2(_11408_),
    .ZN(_11409_));
 CLKBUF_X2 _21098_ (.A(_11340_),
    .Z(_11410_));
 OAI21_X1 _21099_ (.A(_11406_),
    .B1(_11409_),
    .B2(_11410_),
    .ZN(_11411_));
 AND4_X1 _21100_ (.A1(_11392_),
    .A2(_11402_),
    .A3(_11404_),
    .A4(_11411_),
    .ZN(_11412_));
 AND2_X1 _21101_ (.A1(_11316_),
    .A2(_11365_),
    .ZN(_11413_));
 BUF_X2 _21102_ (.A(_11413_),
    .Z(_11414_));
 BUF_X2 _21103_ (.A(_11414_),
    .Z(_11415_));
 INV_X1 _21104_ (.A(_11415_),
    .ZN(_11416_));
 AOI21_X1 _21105_ (.A(_11373_),
    .B1(_11356_),
    .B2(_11408_),
    .ZN(_11417_));
 BUF_X2 _21106_ (.A(_11379_),
    .Z(_11418_));
 AND2_X1 _21107_ (.A1(_11418_),
    .A2(_11320_),
    .ZN(_11419_));
 BUF_X2 _21108_ (.A(_11419_),
    .Z(_11420_));
 NOR2_X1 _21109_ (.A1(_11400_),
    .A2(_11420_),
    .ZN(_11421_));
 AOI21_X1 _21110_ (.A(_11416_),
    .B1(_11417_),
    .B2(_11421_),
    .ZN(_11422_));
 CLKBUF_X2 _21111_ (.A(_11354_),
    .Z(_11423_));
 AND2_X1 _21112_ (.A1(_11423_),
    .A2(_11343_),
    .ZN(_11424_));
 CLKBUF_X2 _21113_ (.A(_11424_),
    .Z(_11425_));
 AND2_X1 _21114_ (.A1(_11365_),
    .A2(_11350_),
    .ZN(_11426_));
 CLKBUF_X2 _21115_ (.A(_11426_),
    .Z(_11427_));
 AND2_X1 _21116_ (.A1(_11425_),
    .A2(_11427_),
    .ZN(_11428_));
 AND2_X1 _21117_ (.A1(_11361_),
    .A2(_11423_),
    .ZN(_11429_));
 AND2_X1 _21118_ (.A1(_11429_),
    .A2(_11426_),
    .ZN(_11430_));
 BUF_X2 _21119_ (.A(_11427_),
    .Z(_11431_));
 AND2_X1 _21120_ (.A1(_11336_),
    .A2(_11431_),
    .ZN(_11432_));
 NOR4_X1 _21121_ (.A1(_11422_),
    .A2(_11428_),
    .A3(_11430_),
    .A4(_11432_),
    .ZN(_11433_));
 BUF_X2 _21122_ (.A(_11366_),
    .Z(_11434_));
 BUF_X2 _21123_ (.A(_11325_),
    .Z(_11435_));
 AND2_X1 _21124_ (.A1(_11395_),
    .A2(_11435_),
    .ZN(_11436_));
 BUF_X2 _21125_ (.A(_11436_),
    .Z(_11437_));
 AND2_X1 _21126_ (.A1(_11434_),
    .A2(_11437_),
    .ZN(_11438_));
 INV_X1 _21127_ (.A(_11438_),
    .ZN(_11439_));
 INV_X1 _21128_ (.A(_11366_),
    .ZN(_11440_));
 INV_X1 _21129_ (.A(_11321_),
    .ZN(_11441_));
 AND2_X1 _21130_ (.A1(_11320_),
    .A2(_11343_),
    .ZN(_11442_));
 INV_X1 _21131_ (.A(_11442_),
    .ZN(_11443_));
 NAND2_X1 _21132_ (.A1(_11441_),
    .A2(_11443_),
    .ZN(_11444_));
 INV_X1 _21133_ (.A(_11444_),
    .ZN(_11445_));
 OAI21_X1 _21134_ (.A(_11439_),
    .B1(_11440_),
    .B2(_11445_),
    .ZN(_11446_));
 OAI21_X1 _21135_ (.A(_11332_),
    .B1(_11388_),
    .B2(_16745_),
    .ZN(_11447_));
 AND3_X1 _21136_ (.A1(_11385_),
    .A2(_11351_),
    .A3(_11332_),
    .ZN(_11448_));
 AND2_X1 _21137_ (.A1(_11447_),
    .A2(_11448_),
    .ZN(_11449_));
 AND2_X2 _21138_ (.A1(_11314_),
    .A2(_11350_),
    .ZN(_11450_));
 AND2_X1 _21139_ (.A1(_11379_),
    .A2(_11354_),
    .ZN(_11451_));
 BUF_X2 _21140_ (.A(_11451_),
    .Z(_11452_));
 OAI21_X1 _21141_ (.A(_11450_),
    .B1(_11452_),
    .B2(_11371_),
    .ZN(_11453_));
 NAND4_X1 _21142_ (.A1(_11314_),
    .A2(_11334_),
    .A3(_11335_),
    .A4(_11351_),
    .ZN(_11454_));
 NAND2_X1 _21143_ (.A1(_11453_),
    .A2(_11454_),
    .ZN(_11455_));
 AND2_X1 _21144_ (.A1(_11423_),
    .A2(_16743_),
    .ZN(_11456_));
 NAND2_X1 _21145_ (.A1(_11434_),
    .A2(_11456_),
    .ZN(_11457_));
 AND2_X1 _21146_ (.A1(_11381_),
    .A2(_11365_),
    .ZN(_11458_));
 CLKBUF_X2 _21147_ (.A(_11458_),
    .Z(_11459_));
 BUF_X2 _21148_ (.A(_11459_),
    .Z(_11460_));
 AND2_X2 _21149_ (.A1(_11320_),
    .A2(_16744_),
    .ZN(_11461_));
 NAND2_X1 _21150_ (.A1(_11460_),
    .A2(_11461_),
    .ZN(_11462_));
 INV_X1 _21151_ (.A(_11459_),
    .ZN(_11463_));
 OAI211_X1 _21152_ (.A(_11457_),
    .B(_11462_),
    .C1(_11359_),
    .C2(_11463_),
    .ZN(_11464_));
 NOR4_X1 _21153_ (.A1(_11446_),
    .A2(_11449_),
    .A3(_11455_),
    .A4(_11464_),
    .ZN(_11465_));
 NAND4_X1 _21154_ (.A1(_11384_),
    .A2(_11412_),
    .A3(_11433_),
    .A4(_11465_),
    .ZN(_11466_));
 AND2_X2 _21155_ (.A1(_11395_),
    .A2(_11319_),
    .ZN(_11467_));
 NAND2_X1 _21156_ (.A1(_11347_),
    .A2(_11467_),
    .ZN(_11468_));
 INV_X1 _21157_ (.A(_11320_),
    .ZN(_11469_));
 OAI22_X1 _21158_ (.A1(_11355_),
    .A2(_11388_),
    .B1(_11469_),
    .B2(_11362_),
    .ZN(_11470_));
 AND2_X1 _21159_ (.A1(_11470_),
    .A2(_11382_),
    .ZN(_11471_));
 BUF_X2 _21160_ (.A(_11360_),
    .Z(_11472_));
 AND2_X1 _21161_ (.A1(_11354_),
    .A2(_16744_),
    .ZN(_11473_));
 AND2_X1 _21162_ (.A1(_11473_),
    .A2(_11426_),
    .ZN(_11474_));
 AOI221_X1 _21163_ (.A(_11471_),
    .B1(_11472_),
    .B2(_11474_),
    .C1(_11420_),
    .C2(_11427_),
    .ZN(_11475_));
 AND2_X1 _21164_ (.A1(_11331_),
    .A2(_11452_),
    .ZN(_11476_));
 AND2_X1 _21165_ (.A1(_11329_),
    .A2(_11349_),
    .ZN(_11477_));
 AND2_X1 _21166_ (.A1(_11477_),
    .A2(_11398_),
    .ZN(_11478_));
 AOI211_X1 _21167_ (.A(_11476_),
    .B(_11478_),
    .C1(_11442_),
    .C2(_11406_),
    .ZN(_11479_));
 AND2_X1 _21168_ (.A1(_11364_),
    .A2(_11385_),
    .ZN(_11480_));
 CLKBUF_X2 _21169_ (.A(_11480_),
    .Z(_11481_));
 BUF_X2 _21170_ (.A(_11481_),
    .Z(_11482_));
 BUF_X2 _21171_ (.A(_11386_),
    .Z(_11483_));
 AOI22_X1 _21172_ (.A1(_11482_),
    .A2(_11425_),
    .B1(_11344_),
    .B2(_11483_),
    .ZN(_11484_));
 AND4_X1 _21173_ (.A1(_11468_),
    .A2(_11475_),
    .A3(_11479_),
    .A4(_11484_),
    .ZN(_11485_));
 AND2_X1 _21174_ (.A1(_11385_),
    .A2(_11350_),
    .ZN(_11486_));
 BUF_X2 _21175_ (.A(_11486_),
    .Z(_11487_));
 BUF_X2 _21176_ (.A(_11487_),
    .Z(_11488_));
 AND2_X1 _21177_ (.A1(_11362_),
    .A2(_11334_),
    .ZN(_11489_));
 NOR3_X1 _21178_ (.A1(_11343_),
    .A2(_11376_),
    .A3(_16746_),
    .ZN(_11490_));
 OAI21_X1 _21179_ (.A(_11488_),
    .B1(_11489_),
    .B2(_11490_),
    .ZN(_11491_));
 AND2_X1 _21180_ (.A1(_11361_),
    .A2(_11320_),
    .ZN(_11492_));
 BUF_X2 _21181_ (.A(_11492_),
    .Z(_11493_));
 NAND2_X1 _21182_ (.A1(_11347_),
    .A2(_11493_),
    .ZN(_11494_));
 AND2_X1 _21183_ (.A1(_11331_),
    .A2(_11321_),
    .ZN(_11495_));
 INV_X1 _21184_ (.A(_11495_),
    .ZN(_11496_));
 BUF_X2 _21185_ (.A(_11450_),
    .Z(_11497_));
 NAND2_X1 _21186_ (.A1(_11398_),
    .A2(_11497_),
    .ZN(_11498_));
 AND2_X1 _21187_ (.A1(_11395_),
    .A2(_11379_),
    .ZN(_11499_));
 NAND2_X1 _21188_ (.A1(_11331_),
    .A2(_11499_),
    .ZN(_11500_));
 AND4_X1 _21189_ (.A1(_11494_),
    .A2(_11496_),
    .A3(_11498_),
    .A4(_11500_),
    .ZN(_11501_));
 NAND2_X1 _21190_ (.A1(_11398_),
    .A2(_11460_),
    .ZN(_11502_));
 NAND2_X1 _21191_ (.A1(_11452_),
    .A2(_11459_),
    .ZN(_11503_));
 NAND2_X1 _21192_ (.A1(_11502_),
    .A2(_11503_),
    .ZN(_11504_));
 NOR2_X1 _21193_ (.A1(_11469_),
    .A2(_11319_),
    .ZN(_11505_));
 AND2_X1 _21194_ (.A1(_11480_),
    .A2(_11505_),
    .ZN(_11506_));
 AND2_X1 _21195_ (.A1(_11388_),
    .A2(_11333_),
    .ZN(_11507_));
 AND2_X1 _21196_ (.A1(_11481_),
    .A2(_11507_),
    .ZN(_11508_));
 AND2_X1 _21197_ (.A1(_11493_),
    .A2(_11459_),
    .ZN(_11509_));
 NOR4_X1 _21198_ (.A1(_11504_),
    .A2(_11506_),
    .A3(_11508_),
    .A4(_11509_),
    .ZN(_11510_));
 BUF_X2 _21199_ (.A(_11499_),
    .Z(_11511_));
 OAI21_X1 _21200_ (.A(_11483_),
    .B1(_11511_),
    .B2(_11370_),
    .ZN(_11512_));
 AND4_X1 _21201_ (.A1(_11491_),
    .A2(_11501_),
    .A3(_11510_),
    .A4(_11512_),
    .ZN(_11513_));
 AND2_X1 _21202_ (.A1(_11371_),
    .A2(_11386_),
    .ZN(_11514_));
 INV_X1 _21203_ (.A(_11514_),
    .ZN(_11515_));
 NAND2_X1 _21204_ (.A1(_11347_),
    .A2(_11437_),
    .ZN(_11516_));
 NAND3_X1 _21205_ (.A1(_11327_),
    .A2(_11351_),
    .A3(_11314_),
    .ZN(_11517_));
 AND2_X1 _21206_ (.A1(_11395_),
    .A2(_16744_),
    .ZN(_11518_));
 NAND2_X1 _21207_ (.A1(_11403_),
    .A2(_11518_),
    .ZN(_11519_));
 NAND4_X1 _21208_ (.A1(_11515_),
    .A2(_11516_),
    .A3(_11517_),
    .A4(_11519_),
    .ZN(_11520_));
 AND2_X1 _21209_ (.A1(_11349_),
    .A2(_11316_),
    .ZN(_11521_));
 CLKBUF_X2 _21210_ (.A(_11521_),
    .Z(_11522_));
 INV_X1 _21211_ (.A(_11522_),
    .ZN(_11523_));
 OAI21_X1 _21212_ (.A(_11389_),
    .B1(_11418_),
    .B2(_11362_),
    .ZN(_11524_));
 BUF_X2 _21213_ (.A(_11473_),
    .Z(_11525_));
 INV_X1 _21214_ (.A(_11525_),
    .ZN(_11526_));
 AOI21_X1 _21215_ (.A(_11523_),
    .B1(_11524_),
    .B2(_11526_),
    .ZN(_11527_));
 AND2_X1 _21216_ (.A1(_11395_),
    .A2(_16743_),
    .ZN(_11528_));
 AND2_X1 _21217_ (.A1(_11405_),
    .A2(_11528_),
    .ZN(_11529_));
 AND2_X1 _21218_ (.A1(_11320_),
    .A2(_16743_),
    .ZN(_11530_));
 AND2_X1 _21219_ (.A1(_11405_),
    .A2(_11530_),
    .ZN(_11531_));
 NOR4_X1 _21220_ (.A1(_11520_),
    .A2(_11527_),
    .A3(_11529_),
    .A4(_11531_),
    .ZN(_11532_));
 AND2_X1 _21221_ (.A1(_11316_),
    .A2(_11385_),
    .ZN(_11533_));
 CLKBUF_X2 _21222_ (.A(_11533_),
    .Z(_11534_));
 AND2_X1 _21223_ (.A1(_11534_),
    .A2(_11461_),
    .ZN(_11535_));
 BUF_X2 _21224_ (.A(_11534_),
    .Z(_11536_));
 AOI21_X1 _21225_ (.A(_11535_),
    .B1(_11346_),
    .B2(_11536_),
    .ZN(_11537_));
 INV_X1 _21226_ (.A(_11499_),
    .ZN(_11538_));
 INV_X1 _21227_ (.A(_11400_),
    .ZN(_11539_));
 NAND2_X2 _21228_ (.A1(_11538_),
    .A2(_11539_),
    .ZN(_11540_));
 OAI21_X1 _21229_ (.A(_11482_),
    .B1(_11540_),
    .B2(_11525_),
    .ZN(_11541_));
 AND2_X1 _21230_ (.A1(_11408_),
    .A2(_11395_),
    .ZN(_11542_));
 NAND3_X1 _21231_ (.A1(_11542_),
    .A2(_11388_),
    .A3(_11536_),
    .ZN(_11543_));
 NOR2_X1 _21232_ (.A1(_11435_),
    .A2(_16745_),
    .ZN(_11544_));
 OAI21_X1 _21233_ (.A(_11488_),
    .B1(_11409_),
    .B2(_11544_),
    .ZN(_11545_));
 AND4_X1 _21234_ (.A1(_11537_),
    .A2(_11541_),
    .A3(_11543_),
    .A4(_11545_),
    .ZN(_11546_));
 NAND4_X1 _21235_ (.A1(_11485_),
    .A2(_11513_),
    .A3(_11532_),
    .A4(_11546_),
    .ZN(_11547_));
 NOR2_X2 _21236_ (.A1(_11466_),
    .A2(_11547_),
    .ZN(_11548_));
 XNOR2_X1 _21237_ (.A(_11312_),
    .B(_11548_),
    .ZN(_11549_));
 INV_X1 _21238_ (.A(_16702_),
    .ZN(_11550_));
 AND2_X1 _21239_ (.A1(_11550_),
    .A2(_16701_),
    .ZN(_11551_));
 NOR2_X2 _21240_ (.A1(_16700_),
    .A2(_16699_),
    .ZN(_11552_));
 AND2_X2 _21241_ (.A1(_11551_),
    .A2(_11552_),
    .ZN(_11553_));
 INV_X2 _21242_ (.A(_16697_),
    .ZN(_11554_));
 NOR2_X2 _21243_ (.A1(_11554_),
    .A2(_16698_),
    .ZN(_11555_));
 NOR2_X2 _21244_ (.A1(_16695_),
    .A2(_16696_),
    .ZN(_11556_));
 AND2_X1 _21245_ (.A1(_11555_),
    .A2(_11556_),
    .ZN(_11557_));
 AND2_X1 _21246_ (.A1(_11553_),
    .A2(_11557_),
    .ZN(_11558_));
 INV_X2 _21247_ (.A(_16696_),
    .ZN(_11559_));
 NOR2_X1 _21248_ (.A1(_11559_),
    .A2(_16695_),
    .ZN(_11560_));
 AND2_X1 _21249_ (.A1(_16698_),
    .A2(_16697_),
    .ZN(_11561_));
 CLKBUF_X2 _21250_ (.A(_11561_),
    .Z(_11562_));
 AND2_X1 _21251_ (.A1(_11560_),
    .A2(_11562_),
    .ZN(_11563_));
 AND2_X2 _21252_ (.A1(_11562_),
    .A2(_11559_),
    .ZN(_11564_));
 OAI21_X1 _21253_ (.A(_11553_),
    .B1(_11563_),
    .B2(_11564_),
    .ZN(_11565_));
 CLKBUF_X2 _21254_ (.A(_11551_),
    .Z(_11566_));
 CLKBUF_X2 _21255_ (.A(_16695_),
    .Z(_11567_));
 INV_X1 _21256_ (.A(_16698_),
    .ZN(_11568_));
 NOR2_X1 _21257_ (.A1(_11568_),
    .A2(_16697_),
    .ZN(_11569_));
 CLKBUF_X2 _21258_ (.A(_11569_),
    .Z(_11570_));
 CLKBUF_X2 _21259_ (.A(_11570_),
    .Z(_11571_));
 CLKBUF_X2 _21260_ (.A(_11552_),
    .Z(_11572_));
 NAND4_X1 _21261_ (.A1(_11566_),
    .A2(_11567_),
    .A3(_11571_),
    .A4(_11572_),
    .ZN(_11573_));
 NAND2_X1 _21262_ (.A1(_11565_),
    .A2(_11573_),
    .ZN(_11574_));
 NOR2_X2 _21263_ (.A1(_16698_),
    .A2(_16697_),
    .ZN(_11575_));
 AND2_X1 _21264_ (.A1(_11575_),
    .A2(_11559_),
    .ZN(_11576_));
 BUF_X2 _21265_ (.A(_11576_),
    .Z(_11577_));
 AOI211_X1 _21266_ (.A(_11558_),
    .B(_11574_),
    .C1(_11553_),
    .C2(_11577_),
    .ZN(_11578_));
 AND2_X1 _21267_ (.A1(_16700_),
    .A2(_16699_),
    .ZN(_11579_));
 AND2_X1 _21268_ (.A1(_11551_),
    .A2(_11579_),
    .ZN(_11580_));
 BUF_X2 _21269_ (.A(_11580_),
    .Z(_11581_));
 INV_X1 _21270_ (.A(_11556_),
    .ZN(_11582_));
 AND2_X2 _21271_ (.A1(_16695_),
    .A2(_16696_),
    .ZN(_11583_));
 NOR3_X1 _21272_ (.A1(_11583_),
    .A2(_11568_),
    .A3(_11554_),
    .ZN(_11584_));
 NAND3_X1 _21273_ (.A1(_11581_),
    .A2(_11582_),
    .A3(_11584_),
    .ZN(_11585_));
 AND2_X1 _21274_ (.A1(_11570_),
    .A2(_11583_),
    .ZN(_11586_));
 CLKBUF_X2 _21275_ (.A(_11586_),
    .Z(_11587_));
 CLKBUF_X2 _21276_ (.A(_11579_),
    .Z(_11588_));
 NAND3_X1 _21277_ (.A1(_11587_),
    .A2(_11588_),
    .A3(_11566_),
    .ZN(_11589_));
 NAND2_X1 _21278_ (.A1(_11585_),
    .A2(_11589_),
    .ZN(_11590_));
 INV_X1 _21279_ (.A(_11580_),
    .ZN(_11591_));
 CLKBUF_X2 _21280_ (.A(_11575_),
    .Z(_11592_));
 AND2_X1 _21281_ (.A1(_11583_),
    .A2(_11592_),
    .ZN(_11593_));
 INV_X1 _21282_ (.A(_11593_),
    .ZN(_11594_));
 INV_X1 _21283_ (.A(_11576_),
    .ZN(_11595_));
 AOI21_X1 _21284_ (.A(_11591_),
    .B1(_11594_),
    .B2(_11595_),
    .ZN(_11596_));
 AND2_X1 _21285_ (.A1(_11555_),
    .A2(_16695_),
    .ZN(_11597_));
 BUF_X2 _21286_ (.A(_11597_),
    .Z(_11598_));
 AOI211_X1 _21287_ (.A(_11590_),
    .B(_11596_),
    .C1(_11581_),
    .C2(_11598_),
    .ZN(_11599_));
 INV_X1 _21288_ (.A(_16699_),
    .ZN(_11600_));
 NOR2_X1 _21289_ (.A1(_11600_),
    .A2(_16700_),
    .ZN(_11601_));
 CLKBUF_X2 _21290_ (.A(_11601_),
    .Z(_11602_));
 AND2_X1 _21291_ (.A1(_11551_),
    .A2(_11602_),
    .ZN(_11603_));
 AND2_X1 _21292_ (.A1(_11555_),
    .A2(_16696_),
    .ZN(_11604_));
 AND2_X1 _21293_ (.A1(_11603_),
    .A2(_11604_),
    .ZN(_11605_));
 INV_X1 _21294_ (.A(_11605_),
    .ZN(_11606_));
 BUF_X2 _21295_ (.A(_11603_),
    .Z(_11607_));
 AND2_X1 _21296_ (.A1(_11570_),
    .A2(_11567_),
    .ZN(_11608_));
 AND2_X1 _21297_ (.A1(_11562_),
    .A2(_11583_),
    .ZN(_11609_));
 OAI21_X1 _21298_ (.A(_11607_),
    .B1(_11608_),
    .B2(_11609_),
    .ZN(_11610_));
 NAND2_X1 _21299_ (.A1(_11603_),
    .A2(_11577_),
    .ZN(_11611_));
 BUF_X2 _21300_ (.A(_11593_),
    .Z(_11612_));
 NAND2_X1 _21301_ (.A1(_11607_),
    .A2(_11612_),
    .ZN(_11613_));
 AND4_X1 _21302_ (.A1(_11606_),
    .A2(_11610_),
    .A3(_11611_),
    .A4(_11613_),
    .ZN(_11614_));
 AND2_X1 _21303_ (.A1(_11600_),
    .A2(_16700_),
    .ZN(_11615_));
 CLKBUF_X2 _21304_ (.A(_11615_),
    .Z(_11616_));
 AND2_X1 _21305_ (.A1(_11551_),
    .A2(_11616_),
    .ZN(_11617_));
 INV_X1 _21306_ (.A(_11617_),
    .ZN(_11618_));
 INV_X1 _21307_ (.A(_11604_),
    .ZN(_11619_));
 CLKBUF_X2 _21308_ (.A(_11555_),
    .Z(_11620_));
 AND2_X1 _21309_ (.A1(_11620_),
    .A2(_11559_),
    .ZN(_11621_));
 CLKBUF_X2 _21310_ (.A(_11621_),
    .Z(_11622_));
 INV_X1 _21311_ (.A(_11622_),
    .ZN(_11623_));
 AOI21_X1 _21312_ (.A(_11618_),
    .B1(_11619_),
    .B2(_11623_),
    .ZN(_11624_));
 INV_X1 _21313_ (.A(_16695_),
    .ZN(_11625_));
 NOR2_X2 _21314_ (.A1(_11625_),
    .A2(_16696_),
    .ZN(_11626_));
 AND2_X1 _21315_ (.A1(_11626_),
    .A2(_11575_),
    .ZN(_11627_));
 INV_X1 _21316_ (.A(_11627_),
    .ZN(_11628_));
 AOI21_X1 _21317_ (.A(_11618_),
    .B1(_11628_),
    .B2(_11594_),
    .ZN(_11629_));
 AND2_X1 _21318_ (.A1(_11617_),
    .A2(_11563_),
    .ZN(_11630_));
 INV_X1 _21319_ (.A(_11570_),
    .ZN(_11631_));
 CLKBUF_X2 _21320_ (.A(_11560_),
    .Z(_11632_));
 NOR2_X1 _21321_ (.A1(_11631_),
    .A2(_11632_),
    .ZN(_11633_));
 AND2_X1 _21322_ (.A1(_11633_),
    .A2(_11617_),
    .ZN(_11634_));
 NOR4_X1 _21323_ (.A1(_11624_),
    .A2(_11629_),
    .A3(_11630_),
    .A4(_11634_),
    .ZN(_11635_));
 AND4_X1 _21324_ (.A1(_11578_),
    .A2(_11599_),
    .A3(_11614_),
    .A4(_11635_),
    .ZN(_11636_));
 NOR2_X2 _21325_ (.A1(_11550_),
    .A2(_16701_),
    .ZN(_11637_));
 AND2_X1 _21326_ (.A1(_11602_),
    .A2(_11637_),
    .ZN(_11638_));
 CLKBUF_X2 _21327_ (.A(_11638_),
    .Z(_11639_));
 NOR3_X2 _21328_ (.A1(_11583_),
    .A2(_16698_),
    .A3(_16697_),
    .ZN(_11640_));
 AND3_X1 _21329_ (.A1(_11639_),
    .A2(_11582_),
    .A3(_11640_),
    .ZN(_11641_));
 CLKBUF_X2 _21330_ (.A(_16696_),
    .Z(_11642_));
 AND2_X1 _21331_ (.A1(_11562_),
    .A2(_11642_),
    .ZN(_11643_));
 BUF_X2 _21332_ (.A(_11643_),
    .Z(_11644_));
 AOI21_X1 _21333_ (.A(_11641_),
    .B1(_11639_),
    .B2(_11644_),
    .ZN(_11645_));
 CLKBUF_X2 _21334_ (.A(_11637_),
    .Z(_11646_));
 AND4_X1 _21335_ (.A1(_11567_),
    .A2(_11571_),
    .A3(_11646_),
    .A4(_11572_),
    .ZN(_11647_));
 INV_X1 _21336_ (.A(_11555_),
    .ZN(_11648_));
 NOR2_X1 _21337_ (.A1(_11648_),
    .A2(_11632_),
    .ZN(_11649_));
 AND2_X1 _21338_ (.A1(_11637_),
    .A2(_11552_),
    .ZN(_11650_));
 NAND2_X1 _21339_ (.A1(_11649_),
    .A2(_11650_),
    .ZN(_11651_));
 INV_X1 _21340_ (.A(_11650_),
    .ZN(_11652_));
 AND2_X1 _21341_ (.A1(_11592_),
    .A2(_11625_),
    .ZN(_11653_));
 INV_X1 _21342_ (.A(_11653_),
    .ZN(_11654_));
 OAI21_X1 _21343_ (.A(_11651_),
    .B1(_11652_),
    .B2(_11654_),
    .ZN(_11655_));
 BUF_X2 _21344_ (.A(_11650_),
    .Z(_11656_));
 NOR3_X1 _21345_ (.A1(_11556_),
    .A2(_11568_),
    .A3(_11554_),
    .ZN(_11657_));
 AOI211_X1 _21346_ (.A(_11647_),
    .B(_11655_),
    .C1(_11656_),
    .C2(_11657_),
    .ZN(_11658_));
 BUF_X2 _21347_ (.A(_11616_),
    .Z(_11659_));
 OAI211_X1 _21348_ (.A(_11646_),
    .B(_11659_),
    .C1(_11609_),
    .C2(_11564_),
    .ZN(_11660_));
 BUF_X2 _21349_ (.A(_11626_),
    .Z(_11661_));
 NAND4_X1 _21350_ (.A1(_11659_),
    .A2(_11571_),
    .A3(_11661_),
    .A4(_11646_),
    .ZN(_11662_));
 NAND2_X1 _21351_ (.A1(_11660_),
    .A2(_11662_),
    .ZN(_11663_));
 AND2_X1 _21352_ (.A1(_11615_),
    .A2(_11637_),
    .ZN(_11664_));
 AND2_X1 _21353_ (.A1(_11664_),
    .A2(_11557_),
    .ZN(_11665_));
 NOR2_X1 _21354_ (.A1(_11663_),
    .A2(_11665_),
    .ZN(_11666_));
 AND2_X2 _21355_ (.A1(_11637_),
    .A2(_11579_),
    .ZN(_11667_));
 INV_X1 _21356_ (.A(_11575_),
    .ZN(_11668_));
 NOR2_X1 _21357_ (.A1(_11668_),
    .A2(_11626_),
    .ZN(_11669_));
 AND2_X1 _21358_ (.A1(_11667_),
    .A2(_11669_),
    .ZN(_11670_));
 INV_X1 _21359_ (.A(_11632_),
    .ZN(_11671_));
 CLKBUF_X2 _21360_ (.A(_11620_),
    .Z(_11672_));
 AND3_X1 _21361_ (.A1(_11667_),
    .A2(_11671_),
    .A3(_11672_),
    .ZN(_11673_));
 AND2_X2 _21362_ (.A1(_11562_),
    .A2(_11556_),
    .ZN(_11674_));
 BUF_X2 _21363_ (.A(_11667_),
    .Z(_11675_));
 AOI211_X1 _21364_ (.A(_11670_),
    .B(_11673_),
    .C1(_11674_),
    .C2(_11675_),
    .ZN(_11676_));
 AND4_X1 _21365_ (.A1(_11645_),
    .A2(_11658_),
    .A3(_11666_),
    .A4(_11676_),
    .ZN(_11677_));
 NOR2_X1 _21366_ (.A1(_16702_),
    .A2(_16701_),
    .ZN(_11678_));
 AND2_X1 _21367_ (.A1(_11601_),
    .A2(_11678_),
    .ZN(_11679_));
 BUF_X2 _21368_ (.A(_11679_),
    .Z(_11680_));
 AND2_X1 _21369_ (.A1(_11626_),
    .A2(_11555_),
    .ZN(_11681_));
 INV_X1 _21370_ (.A(_11681_),
    .ZN(_11682_));
 AND2_X1 _21371_ (.A1(_11560_),
    .A2(_11555_),
    .ZN(_11683_));
 INV_X1 _21372_ (.A(_11683_),
    .ZN(_11684_));
 NAND2_X1 _21373_ (.A1(_11682_),
    .A2(_11684_),
    .ZN(_11685_));
 AND2_X1 _21374_ (.A1(_11575_),
    .A2(_16696_),
    .ZN(_11686_));
 BUF_X2 _21375_ (.A(_11686_),
    .Z(_11687_));
 OAI21_X1 _21376_ (.A(_11680_),
    .B1(_11685_),
    .B2(_11687_),
    .ZN(_11688_));
 AND2_X2 _21377_ (.A1(_11570_),
    .A2(_11556_),
    .ZN(_11689_));
 NAND2_X1 _21378_ (.A1(_11689_),
    .A2(_11680_),
    .ZN(_11690_));
 INV_X1 _21379_ (.A(_11587_),
    .ZN(_11691_));
 INV_X1 _21380_ (.A(_11679_),
    .ZN(_11692_));
 OAI211_X1 _21381_ (.A(_11688_),
    .B(_11690_),
    .C1(_11691_),
    .C2(_11692_),
    .ZN(_11693_));
 AND2_X2 _21382_ (.A1(_11560_),
    .A2(_11575_),
    .ZN(_11694_));
 CLKBUF_X2 _21383_ (.A(_11678_),
    .Z(_11695_));
 AND2_X1 _21384_ (.A1(_11579_),
    .A2(_11695_),
    .ZN(_11696_));
 AND2_X1 _21385_ (.A1(_11694_),
    .A2(_11696_),
    .ZN(_11697_));
 AND2_X1 _21386_ (.A1(_11592_),
    .A2(_16695_),
    .ZN(_11698_));
 AND2_X1 _21387_ (.A1(_11696_),
    .A2(_11698_),
    .ZN(_11699_));
 NOR2_X1 _21388_ (.A1(_11697_),
    .A2(_11699_),
    .ZN(_11700_));
 BUF_X2 _21389_ (.A(_11632_),
    .Z(_11701_));
 BUF_X2 _21390_ (.A(_11672_),
    .Z(_11702_));
 NAND4_X1 _21391_ (.A1(_11701_),
    .A2(_11702_),
    .A3(_11695_),
    .A4(_11588_),
    .ZN(_11703_));
 BUF_X2 _21392_ (.A(_11696_),
    .Z(_11704_));
 CLKBUF_X2 _21393_ (.A(_11562_),
    .Z(_11705_));
 BUF_X2 _21394_ (.A(_11567_),
    .Z(_11706_));
 CLKBUF_X2 _21395_ (.A(_11559_),
    .Z(_11707_));
 OAI211_X1 _21396_ (.A(_11704_),
    .B(_11705_),
    .C1(_11706_),
    .C2(_11707_),
    .ZN(_11708_));
 BUF_X2 _21397_ (.A(_11570_),
    .Z(_11709_));
 BUF_X2 _21398_ (.A(_11556_),
    .Z(_11710_));
 NAND3_X1 _21399_ (.A1(_11704_),
    .A2(_11709_),
    .A3(_11710_),
    .ZN(_11711_));
 NAND4_X1 _21400_ (.A1(_11700_),
    .A2(_11703_),
    .A3(_11708_),
    .A4(_11711_),
    .ZN(_11712_));
 AND2_X2 _21401_ (.A1(_11678_),
    .A2(_11552_),
    .ZN(_11713_));
 CLKBUF_X2 _21402_ (.A(_11713_),
    .Z(_11714_));
 OAI221_X1 _21403_ (.A(_11714_),
    .B1(_11706_),
    .B2(_11642_),
    .C1(_11584_),
    .C2(_11571_),
    .ZN(_11715_));
 OAI211_X1 _21404_ (.A(_11714_),
    .B(_11672_),
    .C1(_11706_),
    .C2(_11642_),
    .ZN(_11716_));
 INV_X1 _21405_ (.A(_11713_),
    .ZN(_11717_));
 INV_X1 _21406_ (.A(_11687_),
    .ZN(_11718_));
 OAI211_X1 _21407_ (.A(_11715_),
    .B(_11716_),
    .C1(_11717_),
    .C2(_11718_),
    .ZN(_11719_));
 NOR2_X1 _21408_ (.A1(_11648_),
    .A2(_11583_),
    .ZN(_11720_));
 AND2_X1 _21409_ (.A1(_11615_),
    .A2(_11678_),
    .ZN(_11721_));
 BUF_X2 _21410_ (.A(_11721_),
    .Z(_11722_));
 NAND3_X1 _21411_ (.A1(_11720_),
    .A2(_11722_),
    .A3(_11582_),
    .ZN(_11723_));
 OAI211_X1 _21412_ (.A(_11695_),
    .B(_11659_),
    .C1(_11674_),
    .C2(_11644_),
    .ZN(_11724_));
 AND2_X1 _21413_ (.A1(_11582_),
    .A2(_11570_),
    .ZN(_11725_));
 NAND2_X1 _21414_ (.A1(_11721_),
    .A2(_11725_),
    .ZN(_11726_));
 NAND2_X1 _21415_ (.A1(_11721_),
    .A2(_11640_),
    .ZN(_11727_));
 NAND4_X1 _21416_ (.A1(_11723_),
    .A2(_11724_),
    .A3(_11726_),
    .A4(_11727_),
    .ZN(_11728_));
 NOR4_X1 _21417_ (.A1(_11693_),
    .A2(_11712_),
    .A3(_11719_),
    .A4(_11728_),
    .ZN(_11729_));
 AND2_X1 _21418_ (.A1(_16702_),
    .A2(_16701_),
    .ZN(_11730_));
 CLKBUF_X2 _21419_ (.A(_11730_),
    .Z(_11731_));
 CLKBUF_X2 _21420_ (.A(_11731_),
    .Z(_11732_));
 NAND4_X1 _21421_ (.A1(_11584_),
    .A2(_11602_),
    .A3(_11732_),
    .A4(_11582_),
    .ZN(_11733_));
 AND2_X1 _21422_ (.A1(_11602_),
    .A2(_11731_),
    .ZN(_11734_));
 BUF_X2 _21423_ (.A(_11734_),
    .Z(_11735_));
 AND2_X1 _21424_ (.A1(_11569_),
    .A2(_11559_),
    .ZN(_11736_));
 BUF_X2 _21425_ (.A(_11736_),
    .Z(_11737_));
 NAND2_X1 _21426_ (.A1(_11735_),
    .A2(_11737_),
    .ZN(_11738_));
 INV_X1 _21427_ (.A(_11734_),
    .ZN(_11739_));
 AND2_X1 _21428_ (.A1(_11569_),
    .A2(_16696_),
    .ZN(_11740_));
 INV_X2 _21429_ (.A(_11740_),
    .ZN(_11741_));
 OAI211_X1 _21430_ (.A(_11733_),
    .B(_11738_),
    .C1(_11739_),
    .C2(_11741_),
    .ZN(_11742_));
 AND2_X1 _21431_ (.A1(_11731_),
    .A2(_11552_),
    .ZN(_11743_));
 NAND3_X1 _21432_ (.A1(_11743_),
    .A2(_11567_),
    .A3(_11571_),
    .ZN(_11744_));
 NAND4_X1 _21433_ (.A1(_11632_),
    .A2(_11731_),
    .A3(_11705_),
    .A4(_11552_),
    .ZN(_11745_));
 INV_X1 _21434_ (.A(_11564_),
    .ZN(_11746_));
 INV_X1 _21435_ (.A(_11743_),
    .ZN(_11747_));
 OAI211_X1 _21436_ (.A(_11744_),
    .B(_11745_),
    .C1(_11746_),
    .C2(_11747_),
    .ZN(_11748_));
 BUF_X2 _21437_ (.A(_11681_),
    .Z(_11749_));
 NAND2_X1 _21438_ (.A1(_11749_),
    .A2(_11734_),
    .ZN(_11750_));
 INV_X1 _21439_ (.A(_11694_),
    .ZN(_11751_));
 OAI21_X1 _21440_ (.A(_11750_),
    .B1(_11739_),
    .B2(_11751_),
    .ZN(_11752_));
 AND4_X1 _21441_ (.A1(_11731_),
    .A2(_11632_),
    .A3(_11592_),
    .A4(_11552_),
    .ZN(_11753_));
 NOR4_X1 _21442_ (.A1(_11742_),
    .A2(_11748_),
    .A3(_11752_),
    .A4(_11753_),
    .ZN(_11754_));
 AND2_X1 _21443_ (.A1(_11615_),
    .A2(_11730_),
    .ZN(_11755_));
 BUF_X2 _21444_ (.A(_11755_),
    .Z(_11756_));
 AND2_X2 _21445_ (.A1(_11575_),
    .A2(_11556_),
    .ZN(_11757_));
 INV_X1 _21446_ (.A(_11757_),
    .ZN(_11758_));
 NAND2_X1 _21447_ (.A1(_11594_),
    .A2(_11758_),
    .ZN(_11759_));
 OAI21_X1 _21448_ (.A(_11756_),
    .B1(_11759_),
    .B2(_11622_),
    .ZN(_11760_));
 NOR2_X1 _21449_ (.A1(_11631_),
    .A2(_11661_),
    .ZN(_11761_));
 AND2_X1 _21450_ (.A1(_11562_),
    .A2(_11567_),
    .ZN(_11762_));
 OAI21_X1 _21451_ (.A(_11756_),
    .B1(_11761_),
    .B2(_11762_),
    .ZN(_11763_));
 AND2_X2 _21452_ (.A1(_11730_),
    .A2(_11579_),
    .ZN(_11764_));
 AND2_X1 _21453_ (.A1(_11557_),
    .A2(_11764_),
    .ZN(_11765_));
 INV_X1 _21454_ (.A(_11765_),
    .ZN(_11766_));
 BUF_X2 _21455_ (.A(_11764_),
    .Z(_11767_));
 BUF_X2 _21456_ (.A(_11740_),
    .Z(_11768_));
 OAI21_X1 _21457_ (.A(_11767_),
    .B1(_11737_),
    .B2(_11768_),
    .ZN(_11769_));
 OAI211_X1 _21458_ (.A(_11767_),
    .B(_11592_),
    .C1(_11567_),
    .C2(_11642_),
    .ZN(_11770_));
 NAND3_X1 _21459_ (.A1(_11764_),
    .A2(_11632_),
    .A3(_11705_),
    .ZN(_11771_));
 AND4_X1 _21460_ (.A1(_11766_),
    .A2(_11769_),
    .A3(_11770_),
    .A4(_11771_),
    .ZN(_11772_));
 AND4_X1 _21461_ (.A1(_11754_),
    .A2(_11760_),
    .A3(_11763_),
    .A4(_11772_),
    .ZN(_11773_));
 NAND4_X1 _21462_ (.A1(_11636_),
    .A2(_11677_),
    .A3(_11729_),
    .A4(_11773_),
    .ZN(_11774_));
 AND2_X2 _21463_ (.A1(_11714_),
    .A2(_11757_),
    .ZN(_11775_));
 NOR2_X2 _21464_ (.A1(_11774_),
    .A2(_11775_),
    .ZN(_11776_));
 AND2_X1 _21465_ (.A1(_11569_),
    .A2(_11626_),
    .ZN(_11777_));
 INV_X1 _21466_ (.A(_11777_),
    .ZN(_11778_));
 AND2_X1 _21467_ (.A1(_11569_),
    .A2(_11560_),
    .ZN(_11779_));
 INV_X1 _21468_ (.A(_11779_),
    .ZN(_11780_));
 NAND2_X1 _21469_ (.A1(_11778_),
    .A2(_11780_),
    .ZN(_11781_));
 AND2_X1 _21470_ (.A1(_11781_),
    .A2(_11638_),
    .ZN(_11782_));
 INV_X1 _21471_ (.A(_11638_),
    .ZN(_11783_));
 INV_X1 _21472_ (.A(_11698_),
    .ZN(_11784_));
 AOI21_X1 _21473_ (.A(_11783_),
    .B1(_11784_),
    .B2(_11619_),
    .ZN(_11785_));
 INV_X1 _21474_ (.A(_11562_),
    .ZN(_11786_));
 NOR2_X1 _21475_ (.A1(_11786_),
    .A2(_11632_),
    .ZN(_11787_));
 INV_X2 _21476_ (.A(_11626_),
    .ZN(_11788_));
 AND3_X1 _21477_ (.A1(_11639_),
    .A2(_11787_),
    .A3(_11788_),
    .ZN(_11789_));
 NOR3_X1 _21478_ (.A1(_11782_),
    .A2(_11785_),
    .A3(_11789_),
    .ZN(_11790_));
 AND2_X1 _21479_ (.A1(_11683_),
    .A2(_11734_),
    .ZN(_11791_));
 AND2_X1 _21480_ (.A1(_11734_),
    .A2(_11694_),
    .ZN(_11792_));
 NOR2_X1 _21481_ (.A1(_11791_),
    .A2(_11792_),
    .ZN(_11793_));
 AND2_X1 _21482_ (.A1(_11734_),
    .A2(_11586_),
    .ZN(_11794_));
 INV_X1 _21483_ (.A(_11794_),
    .ZN(_11795_));
 INV_X1 _21484_ (.A(_11787_),
    .ZN(_11796_));
 OAI211_X1 _21485_ (.A(_11793_),
    .B(_11795_),
    .C1(_11739_),
    .C2(_11796_),
    .ZN(_11797_));
 OAI21_X1 _21486_ (.A(_11764_),
    .B1(_11621_),
    .B2(_11640_),
    .ZN(_11798_));
 AND2_X1 _21487_ (.A1(_11562_),
    .A2(_11625_),
    .ZN(_11799_));
 NAND2_X1 _21488_ (.A1(_11767_),
    .A2(_11799_),
    .ZN(_11800_));
 INV_X1 _21489_ (.A(_11764_),
    .ZN(_11801_));
 OAI211_X1 _21490_ (.A(_11798_),
    .B(_11800_),
    .C1(_11778_),
    .C2(_11801_),
    .ZN(_11802_));
 OAI211_X1 _21491_ (.A(_11755_),
    .B(_11788_),
    .C1(_11787_),
    .C2(_11570_),
    .ZN(_11803_));
 NAND2_X1 _21492_ (.A1(_11756_),
    .A2(_11604_),
    .ZN(_11804_));
 OAI21_X1 _21493_ (.A(_11755_),
    .B1(_11694_),
    .B2(_11576_),
    .ZN(_11805_));
 NAND3_X1 _21494_ (.A1(_11749_),
    .A2(_11731_),
    .A3(_11616_),
    .ZN(_11806_));
 NAND4_X1 _21495_ (.A1(_11803_),
    .A2(_11804_),
    .A3(_11805_),
    .A4(_11806_),
    .ZN(_11807_));
 OAI211_X1 _21496_ (.A(_11743_),
    .B(_11562_),
    .C1(_11567_),
    .C2(_11642_),
    .ZN(_11808_));
 NOR3_X1 _21497_ (.A1(_11710_),
    .A2(_16698_),
    .A3(_11554_),
    .ZN(_11809_));
 OAI21_X1 _21498_ (.A(_11743_),
    .B1(_11809_),
    .B2(_11757_),
    .ZN(_11810_));
 INV_X2 _21499_ (.A(_11736_),
    .ZN(_11811_));
 OAI211_X1 _21500_ (.A(_11808_),
    .B(_11810_),
    .C1(_11811_),
    .C2(_11747_),
    .ZN(_11812_));
 NOR4_X1 _21501_ (.A1(_11797_),
    .A2(_11802_),
    .A3(_11807_),
    .A4(_11812_),
    .ZN(_11813_));
 AND4_X1 _21502_ (.A1(_11661_),
    .A2(_11620_),
    .A3(_11637_),
    .A4(_11552_),
    .ZN(_11814_));
 AND2_X1 _21503_ (.A1(_11737_),
    .A2(_11650_),
    .ZN(_11815_));
 AOI211_X1 _21504_ (.A(_11814_),
    .B(_11815_),
    .C1(_11656_),
    .C2(_11759_),
    .ZN(_11816_));
 NOR2_X1 _21505_ (.A1(_11563_),
    .A2(_11768_),
    .ZN(_11817_));
 INV_X1 _21506_ (.A(_11667_),
    .ZN(_11818_));
 NOR2_X1 _21507_ (.A1(_11817_),
    .A2(_11818_),
    .ZN(_11819_));
 INV_X1 _21508_ (.A(_11819_),
    .ZN(_11820_));
 CLKBUF_X2 _21509_ (.A(_11664_),
    .Z(_11821_));
 AND2_X1 _21510_ (.A1(_11821_),
    .A2(_11757_),
    .ZN(_11822_));
 INV_X1 _21511_ (.A(_11822_),
    .ZN(_11823_));
 CLKBUF_X2 _21512_ (.A(_11625_),
    .Z(_11824_));
 OAI221_X1 _21513_ (.A(_11821_),
    .B1(_11824_),
    .B2(_11559_),
    .C1(_11571_),
    .C2(_11705_),
    .ZN(_11825_));
 OAI21_X1 _21514_ (.A(_11667_),
    .B1(_11649_),
    .B2(_11577_),
    .ZN(_11826_));
 AND4_X1 _21515_ (.A1(_11820_),
    .A2(_11823_),
    .A3(_11825_),
    .A4(_11826_),
    .ZN(_11827_));
 AND4_X1 _21516_ (.A1(_11790_),
    .A2(_11813_),
    .A3(_11816_),
    .A4(_11827_),
    .ZN(_11828_));
 AND2_X1 _21517_ (.A1(_11580_),
    .A2(_11736_),
    .ZN(_11829_));
 AND2_X1 _21518_ (.A1(_11580_),
    .A2(_11779_),
    .ZN(_11830_));
 AND2_X1 _21519_ (.A1(_11580_),
    .A2(_11657_),
    .ZN(_11831_));
 OR3_X1 _21520_ (.A1(_11829_),
    .A2(_11830_),
    .A3(_11831_),
    .ZN(_11832_));
 AND2_X1 _21521_ (.A1(_11555_),
    .A2(_11583_),
    .ZN(_11833_));
 NAND2_X1 _21522_ (.A1(_11581_),
    .A2(_11833_),
    .ZN(_11834_));
 NAND2_X1 _21523_ (.A1(_11580_),
    .A2(_11621_),
    .ZN(_11835_));
 OAI211_X1 _21524_ (.A(_11834_),
    .B(_11835_),
    .C1(_11591_),
    .C2(_11784_),
    .ZN(_11836_));
 NAND2_X1 _21525_ (.A1(_11617_),
    .A2(_11687_),
    .ZN(_11837_));
 NAND2_X1 _21526_ (.A1(_11617_),
    .A2(_11833_),
    .ZN(_11838_));
 OAI211_X1 _21527_ (.A(_11837_),
    .B(_11838_),
    .C1(_11618_),
    .C2(_11595_),
    .ZN(_11839_));
 INV_X1 _21528_ (.A(_11643_),
    .ZN(_11840_));
 AOI21_X1 _21529_ (.A(_11618_),
    .B1(_11778_),
    .B2(_11840_),
    .ZN(_11841_));
 NOR4_X1 _21530_ (.A1(_11832_),
    .A2(_11836_),
    .A3(_11839_),
    .A4(_11841_),
    .ZN(_11842_));
 INV_X1 _21531_ (.A(_11603_),
    .ZN(_11843_));
 INV_X1 _21532_ (.A(_11781_),
    .ZN(_11844_));
 INV_X1 _21533_ (.A(_11609_),
    .ZN(_11845_));
 AOI21_X1 _21534_ (.A(_11843_),
    .B1(_11844_),
    .B2(_11845_),
    .ZN(_11846_));
 INV_X2 _21535_ (.A(_11553_),
    .ZN(_11847_));
 INV_X1 _21536_ (.A(_11833_),
    .ZN(_11848_));
 AOI21_X1 _21537_ (.A(_11847_),
    .B1(_11628_),
    .B2(_11848_),
    .ZN(_11849_));
 INV_X1 _21538_ (.A(_11762_),
    .ZN(_11850_));
 AOI21_X1 _21539_ (.A(_11847_),
    .B1(_11741_),
    .B2(_11850_),
    .ZN(_11851_));
 OAI21_X1 _21540_ (.A(_11603_),
    .B1(_11749_),
    .B2(_11683_),
    .ZN(_11852_));
 OAI21_X1 _21541_ (.A(_11852_),
    .B1(_11784_),
    .B2(_11843_),
    .ZN(_11853_));
 NOR4_X1 _21542_ (.A1(_11846_),
    .A2(_11849_),
    .A3(_11851_),
    .A4(_11853_),
    .ZN(_11854_));
 NAND3_X1 _21543_ (.A1(_11649_),
    .A2(_11788_),
    .A3(_11680_),
    .ZN(_11855_));
 NAND3_X1 _21544_ (.A1(_11576_),
    .A2(_11602_),
    .A3(_11695_),
    .ZN(_11856_));
 OAI211_X1 _21545_ (.A(_11855_),
    .B(_11856_),
    .C1(_11751_),
    .C2(_11692_),
    .ZN(_11857_));
 NAND4_X1 _21546_ (.A1(_11713_),
    .A2(_11671_),
    .A3(_11788_),
    .A4(_11620_),
    .ZN(_11858_));
 NAND2_X1 _21547_ (.A1(_11564_),
    .A2(_11713_),
    .ZN(_11859_));
 INV_X1 _21548_ (.A(_11563_),
    .ZN(_11860_));
 OAI211_X1 _21549_ (.A(_11858_),
    .B(_11859_),
    .C1(_11860_),
    .C2(_11717_),
    .ZN(_11861_));
 AOI21_X1 _21550_ (.A(_11692_),
    .B1(_11811_),
    .B2(_11741_),
    .ZN(_11862_));
 AOI21_X1 _21551_ (.A(_11692_),
    .B1(_11845_),
    .B2(_11746_),
    .ZN(_11863_));
 NOR4_X1 _21552_ (.A1(_11857_),
    .A2(_11861_),
    .A3(_11862_),
    .A4(_11863_),
    .ZN(_11864_));
 AND2_X1 _21553_ (.A1(_11721_),
    .A2(_11604_),
    .ZN(_11865_));
 INV_X1 _21554_ (.A(_11865_),
    .ZN(_11866_));
 AND2_X1 _21555_ (.A1(_11626_),
    .A2(_11561_),
    .ZN(_11867_));
 AND3_X1 _21556_ (.A1(_11867_),
    .A2(_11695_),
    .A3(_11616_),
    .ZN(_11868_));
 INV_X1 _21557_ (.A(_11868_),
    .ZN(_11869_));
 NAND4_X1 _21558_ (.A1(_11866_),
    .A2(_11869_),
    .A3(_11726_),
    .A4(_11727_),
    .ZN(_11870_));
 AND2_X1 _21559_ (.A1(_11598_),
    .A2(_11696_),
    .ZN(_11871_));
 INV_X1 _21560_ (.A(_11696_),
    .ZN(_11872_));
 INV_X1 _21561_ (.A(_11799_),
    .ZN(_11873_));
 AOI21_X1 _21562_ (.A(_11872_),
    .B1(_11741_),
    .B2(_11873_),
    .ZN(_11874_));
 NOR4_X1 _21563_ (.A1(_11870_),
    .A2(_11699_),
    .A3(_11871_),
    .A4(_11874_),
    .ZN(_11875_));
 AND4_X1 _21564_ (.A1(_11842_),
    .A2(_11854_),
    .A3(_11864_),
    .A4(_11875_),
    .ZN(_11876_));
 AND2_X2 _21565_ (.A1(_11828_),
    .A2(_11876_),
    .ZN(_11877_));
 XOR2_X2 _21566_ (.A(_11776_),
    .B(_11877_),
    .Z(_11878_));
 XNOR2_X1 _21567_ (.A(_11549_),
    .B(_11878_),
    .ZN(_11879_));
 INV_X1 _21568_ (.A(_16785_),
    .ZN(_11880_));
 NOR2_X2 _21569_ (.A1(_11880_),
    .A2(_16786_),
    .ZN(_11881_));
 AND2_X1 _21570_ (.A1(_11881_),
    .A2(_16784_),
    .ZN(_11882_));
 INV_X1 _21571_ (.A(_16788_),
    .ZN(_11883_));
 NOR2_X1 _21572_ (.A1(_11883_),
    .A2(_16787_),
    .ZN(_11884_));
 AND2_X1 _21573_ (.A1(_16790_),
    .A2(_16789_),
    .ZN(_11885_));
 AND2_X1 _21574_ (.A1(_11884_),
    .A2(_11885_),
    .ZN(_11886_));
 CLKBUF_X2 _21575_ (.A(_11886_),
    .Z(_11887_));
 AND2_X1 _21576_ (.A1(_11882_),
    .A2(_11887_),
    .ZN(_11888_));
 INV_X1 _21577_ (.A(_16784_),
    .ZN(_11889_));
 BUF_X2 _21578_ (.A(_16783_),
    .Z(_11890_));
 NOR2_X2 _21579_ (.A1(_11889_),
    .A2(_11890_),
    .ZN(_11891_));
 NOR2_X1 _21580_ (.A1(_16786_),
    .A2(_16785_),
    .ZN(_11892_));
 CLKBUF_X2 _21581_ (.A(_11892_),
    .Z(_11893_));
 AND2_X2 _21582_ (.A1(_11891_),
    .A2(_11893_),
    .ZN(_11894_));
 AND2_X1 _21583_ (.A1(_11894_),
    .A2(_11887_),
    .ZN(_11895_));
 INV_X1 _21584_ (.A(_16783_),
    .ZN(_11896_));
 NOR2_X1 _21585_ (.A1(_11896_),
    .A2(_16784_),
    .ZN(_11897_));
 AND2_X2 _21586_ (.A1(_11897_),
    .A2(_11881_),
    .ZN(_11898_));
 AND2_X1 _21587_ (.A1(_11898_),
    .A2(_11887_),
    .ZN(_11899_));
 AND2_X2 _21588_ (.A1(_11892_),
    .A2(_11889_),
    .ZN(_11900_));
 AND2_X1 _21589_ (.A1(_11886_),
    .A2(_11900_),
    .ZN(_11901_));
 OR4_X1 _21590_ (.A1(_11888_),
    .A2(_11895_),
    .A3(_11899_),
    .A4(_11901_),
    .ZN(_11902_));
 AND2_X1 _21591_ (.A1(_16786_),
    .A2(_16785_),
    .ZN(_11903_));
 CLKBUF_X2 _21592_ (.A(_11903_),
    .Z(_11904_));
 NOR2_X1 _21593_ (.A1(_16783_),
    .A2(_16784_),
    .ZN(_11905_));
 CLKBUF_X2 _21594_ (.A(_11905_),
    .Z(_11906_));
 AND2_X1 _21595_ (.A1(_11904_),
    .A2(_11906_),
    .ZN(_11907_));
 AND2_X1 _21596_ (.A1(_11887_),
    .A2(_11907_),
    .ZN(_11908_));
 AND2_X2 _21597_ (.A1(_11890_),
    .A2(_16784_),
    .ZN(_11909_));
 AND2_X1 _21598_ (.A1(_11909_),
    .A2(_11903_),
    .ZN(_11910_));
 CLKBUF_X2 _21599_ (.A(_11884_),
    .Z(_11911_));
 BUF_X2 _21600_ (.A(_11885_),
    .Z(_11912_));
 AND3_X1 _21601_ (.A1(_11910_),
    .A2(_11911_),
    .A3(_11912_),
    .ZN(_11913_));
 NOR2_X1 _21602_ (.A1(_11908_),
    .A2(_11913_),
    .ZN(_11914_));
 INV_X1 _21603_ (.A(_11914_),
    .ZN(_11915_));
 INV_X1 _21604_ (.A(_16786_),
    .ZN(_11916_));
 NOR2_X1 _21605_ (.A1(_11916_),
    .A2(_16785_),
    .ZN(_11917_));
 CLKBUF_X2 _21606_ (.A(_11917_),
    .Z(_11918_));
 BUF_X2 _21607_ (.A(_11909_),
    .Z(_11919_));
 CLKBUF_X2 _21608_ (.A(_11891_),
    .Z(_11920_));
 OAI211_X1 _21609_ (.A(_11887_),
    .B(_11918_),
    .C1(_11919_),
    .C2(_11920_),
    .ZN(_11921_));
 NAND4_X1 _21610_ (.A1(_11911_),
    .A2(_11918_),
    .A3(_11906_),
    .A4(_11912_),
    .ZN(_11922_));
 NAND2_X1 _21611_ (.A1(_11921_),
    .A2(_11922_),
    .ZN(_11923_));
 AND2_X1 _21612_ (.A1(_16788_),
    .A2(_16787_),
    .ZN(_11924_));
 AND2_X1 _21613_ (.A1(_11912_),
    .A2(_11924_),
    .ZN(_11925_));
 BUF_X2 _21614_ (.A(_11925_),
    .Z(_11926_));
 CLKBUF_X2 _21615_ (.A(_11897_),
    .Z(_11927_));
 AND2_X1 _21616_ (.A1(_11917_),
    .A2(_11927_),
    .ZN(_11928_));
 BUF_X2 _21617_ (.A(_11928_),
    .Z(_11929_));
 AND2_X1 _21618_ (.A1(_11904_),
    .A2(_11896_),
    .ZN(_11930_));
 OAI21_X1 _21619_ (.A(_11926_),
    .B1(_11929_),
    .B2(_11930_),
    .ZN(_11931_));
 CLKBUF_X2 _21620_ (.A(_11896_),
    .Z(_11932_));
 CLKBUF_X2 _21621_ (.A(_11889_),
    .Z(_11933_));
 OAI211_X1 _21622_ (.A(_11926_),
    .B(_11893_),
    .C1(_11932_),
    .C2(_11933_),
    .ZN(_11934_));
 INV_X1 _21623_ (.A(_11926_),
    .ZN(_11935_));
 AND2_X1 _21624_ (.A1(_11881_),
    .A2(_11889_),
    .ZN(_11936_));
 BUF_X2 _21625_ (.A(_11936_),
    .Z(_11937_));
 INV_X1 _21626_ (.A(_11937_),
    .ZN(_11938_));
 OAI211_X1 _21627_ (.A(_11931_),
    .B(_11934_),
    .C1(_11935_),
    .C2(_11938_),
    .ZN(_11939_));
 NOR4_X1 _21628_ (.A1(_11902_),
    .A2(_11915_),
    .A3(_11923_),
    .A4(_11939_),
    .ZN(_11940_));
 NOR2_X2 _21629_ (.A1(_16788_),
    .A2(_16787_),
    .ZN(_11941_));
 AND2_X2 _21630_ (.A1(_11885_),
    .A2(_11941_),
    .ZN(_11942_));
 BUF_X2 _21631_ (.A(_11942_),
    .Z(_11943_));
 BUF_X2 _21632_ (.A(_11881_),
    .Z(_11944_));
 BUF_X2 _21633_ (.A(_11890_),
    .Z(_11945_));
 CLKBUF_X2 _21634_ (.A(_16784_),
    .Z(_11946_));
 OAI211_X1 _21635_ (.A(_11943_),
    .B(_11944_),
    .C1(_11945_),
    .C2(_11946_),
    .ZN(_11947_));
 AND2_X1 _21636_ (.A1(_11903_),
    .A2(_16784_),
    .ZN(_11948_));
 AND2_X1 _21637_ (.A1(_11942_),
    .A2(_11948_),
    .ZN(_11949_));
 AND2_X1 _21638_ (.A1(_11917_),
    .A2(_11889_),
    .ZN(_11950_));
 AND2_X1 _21639_ (.A1(_11950_),
    .A2(_11942_),
    .ZN(_11951_));
 AND2_X1 _21640_ (.A1(_11927_),
    .A2(_11904_),
    .ZN(_11952_));
 BUF_X2 _21641_ (.A(_11952_),
    .Z(_11953_));
 AOI211_X1 _21642_ (.A(_11949_),
    .B(_11951_),
    .C1(_11953_),
    .C2(_11942_),
    .ZN(_11954_));
 BUF_X2 _21643_ (.A(_11893_),
    .Z(_11955_));
 NAND4_X1 _21644_ (.A1(_11912_),
    .A2(_11906_),
    .A3(_11955_),
    .A4(_11941_),
    .ZN(_11956_));
 AND2_X2 _21645_ (.A1(_11883_),
    .A2(_16787_),
    .ZN(_11957_));
 AND2_X1 _21646_ (.A1(_11957_),
    .A2(_11885_),
    .ZN(_11958_));
 BUF_X2 _21647_ (.A(_11958_),
    .Z(_11959_));
 NAND2_X1 _21648_ (.A1(_11959_),
    .A2(_11894_),
    .ZN(_11960_));
 OAI211_X1 _21649_ (.A(_11959_),
    .B(_11904_),
    .C1(_11890_),
    .C2(_11933_),
    .ZN(_11961_));
 AND2_X1 _21650_ (.A1(_11891_),
    .A2(_11881_),
    .ZN(_11962_));
 NAND2_X1 _21651_ (.A1(_11959_),
    .A2(_11962_),
    .ZN(_11963_));
 AND2_X2 _21652_ (.A1(_11917_),
    .A2(_11909_),
    .ZN(_11964_));
 NAND2_X1 _21653_ (.A1(_11959_),
    .A2(_11964_),
    .ZN(_11965_));
 AND4_X1 _21654_ (.A1(_11960_),
    .A2(_11961_),
    .A3(_11963_),
    .A4(_11965_),
    .ZN(_11966_));
 AND4_X1 _21655_ (.A1(_11947_),
    .A2(_11954_),
    .A3(_11956_),
    .A4(_11966_),
    .ZN(_11967_));
 INV_X1 _21656_ (.A(_11905_),
    .ZN(_11968_));
 NAND2_X1 _21657_ (.A1(_11968_),
    .A2(_11918_),
    .ZN(_11969_));
 NOR2_X1 _21658_ (.A1(_11969_),
    .A2(_11909_),
    .ZN(_11970_));
 INV_X1 _21659_ (.A(_16789_),
    .ZN(_11971_));
 AND2_X1 _21660_ (.A1(_11971_),
    .A2(_16790_),
    .ZN(_11972_));
 AND2_X1 _21661_ (.A1(_11972_),
    .A2(_11957_),
    .ZN(_11973_));
 CLKBUF_X2 _21662_ (.A(_11973_),
    .Z(_11974_));
 AND2_X1 _21663_ (.A1(_11970_),
    .A2(_11974_),
    .ZN(_11975_));
 INV_X1 _21664_ (.A(_11975_),
    .ZN(_11976_));
 BUF_X2 _21665_ (.A(_11957_),
    .Z(_11977_));
 CLKBUF_X2 _21666_ (.A(_11972_),
    .Z(_11978_));
 BUF_X2 _21667_ (.A(_11978_),
    .Z(_11979_));
 BUF_X2 _21668_ (.A(_11910_),
    .Z(_11980_));
 OAI211_X1 _21669_ (.A(_11977_),
    .B(_11979_),
    .C1(_11980_),
    .C2(_11907_),
    .ZN(_11981_));
 NAND2_X1 _21670_ (.A1(_11976_),
    .A2(_11981_),
    .ZN(_11982_));
 AND2_X1 _21671_ (.A1(_11978_),
    .A2(_11941_),
    .ZN(_11983_));
 INV_X1 _21672_ (.A(_11983_),
    .ZN(_11984_));
 AND2_X1 _21673_ (.A1(_11909_),
    .A2(_11892_),
    .ZN(_11985_));
 INV_X1 _21674_ (.A(_11985_),
    .ZN(_11986_));
 AND2_X1 _21675_ (.A1(_11905_),
    .A2(_11893_),
    .ZN(_11987_));
 INV_X1 _21676_ (.A(_11987_),
    .ZN(_11988_));
 NAND2_X1 _21677_ (.A1(_11986_),
    .A2(_11988_),
    .ZN(_11989_));
 INV_X1 _21678_ (.A(_11989_),
    .ZN(_11990_));
 INV_X1 _21679_ (.A(_11898_),
    .ZN(_11991_));
 AOI21_X1 _21680_ (.A(_11984_),
    .B1(_11990_),
    .B2(_11991_),
    .ZN(_11992_));
 CLKBUF_X2 _21681_ (.A(_11983_),
    .Z(_11993_));
 CLKBUF_X2 _21682_ (.A(_11950_),
    .Z(_11994_));
 AND2_X1 _21683_ (.A1(_11993_),
    .A2(_11994_),
    .ZN(_11995_));
 NAND4_X1 _21684_ (.A1(_11978_),
    .A2(_11957_),
    .A3(_11944_),
    .A4(_11946_),
    .ZN(_11996_));
 NAND4_X1 _21685_ (.A1(_11977_),
    .A2(_11978_),
    .A3(_11945_),
    .A4(_11893_),
    .ZN(_11997_));
 NAND2_X1 _21686_ (.A1(_11996_),
    .A2(_11997_),
    .ZN(_11998_));
 NOR4_X1 _21687_ (.A1(_11982_),
    .A2(_11992_),
    .A3(_11995_),
    .A4(_11998_),
    .ZN(_11999_));
 AND2_X2 _21688_ (.A1(_11978_),
    .A2(_11924_),
    .ZN(_12000_));
 AND2_X1 _21689_ (.A1(_11917_),
    .A2(_16784_),
    .ZN(_12001_));
 AND2_X1 _21690_ (.A1(_12000_),
    .A2(_12001_),
    .ZN(_12002_));
 AND2_X2 _21691_ (.A1(_11891_),
    .A2(_11904_),
    .ZN(_12003_));
 AND2_X1 _21692_ (.A1(_12000_),
    .A2(_12003_),
    .ZN(_12004_));
 NOR2_X1 _21693_ (.A1(_12002_),
    .A2(_12004_),
    .ZN(_12005_));
 AND2_X1 _21694_ (.A1(_11978_),
    .A2(_11911_),
    .ZN(_12006_));
 AND2_X1 _21695_ (.A1(_12006_),
    .A2(_11987_),
    .ZN(_12007_));
 INV_X1 _21696_ (.A(_12007_),
    .ZN(_12008_));
 CLKBUF_X2 _21697_ (.A(_12006_),
    .Z(_12009_));
 CLKBUF_X2 _21698_ (.A(_11918_),
    .Z(_12010_));
 CLKBUF_X2 _21699_ (.A(_11904_),
    .Z(_12011_));
 OAI221_X1 _21700_ (.A(_12009_),
    .B1(_11932_),
    .B2(_11933_),
    .C1(_12010_),
    .C2(_12011_),
    .ZN(_12012_));
 INV_X1 _21701_ (.A(_11881_),
    .ZN(_12013_));
 NOR2_X1 _21702_ (.A1(_12013_),
    .A2(_11891_),
    .ZN(_12014_));
 OAI21_X1 _21703_ (.A(_12000_),
    .B1(_12014_),
    .B2(_11900_),
    .ZN(_12015_));
 AND4_X1 _21704_ (.A1(_12005_),
    .A2(_12008_),
    .A3(_12012_),
    .A4(_12015_),
    .ZN(_12016_));
 NAND4_X1 _21705_ (.A1(_11940_),
    .A2(_11967_),
    .A3(_11999_),
    .A4(_12016_),
    .ZN(_12017_));
 NOR2_X2 _21706_ (.A1(_16790_),
    .A2(_16789_),
    .ZN(_12018_));
 AND2_X2 _21707_ (.A1(_11957_),
    .A2(_12018_),
    .ZN(_12019_));
 AND2_X1 _21708_ (.A1(_12019_),
    .A2(_12001_),
    .ZN(_12020_));
 INV_X1 _21709_ (.A(_12020_),
    .ZN(_12021_));
 BUF_X2 _21710_ (.A(_12019_),
    .Z(_12022_));
 AND2_X1 _21711_ (.A1(_11904_),
    .A2(_11933_),
    .ZN(_12023_));
 CLKBUF_X2 _21712_ (.A(_12023_),
    .Z(_12024_));
 NAND2_X1 _21713_ (.A1(_12022_),
    .A2(_12024_),
    .ZN(_12025_));
 NAND2_X1 _21714_ (.A1(_12019_),
    .A2(_11980_),
    .ZN(_12026_));
 AND2_X1 _21715_ (.A1(_11918_),
    .A2(_11906_),
    .ZN(_12027_));
 OAI21_X1 _21716_ (.A(_12019_),
    .B1(_11929_),
    .B2(_12027_),
    .ZN(_12028_));
 NAND4_X1 _21717_ (.A1(_12021_),
    .A2(_12025_),
    .A3(_12026_),
    .A4(_12028_),
    .ZN(_12029_));
 AND2_X2 _21718_ (.A1(_12018_),
    .A2(_11941_),
    .ZN(_12030_));
 AND2_X1 _21719_ (.A1(_12003_),
    .A2(_12030_),
    .ZN(_12031_));
 INV_X1 _21720_ (.A(_12031_),
    .ZN(_12032_));
 AND2_X2 _21721_ (.A1(_11881_),
    .A2(_11909_),
    .ZN(_12033_));
 AND2_X2 _21722_ (.A1(_11881_),
    .A2(_11906_),
    .ZN(_12034_));
 OAI21_X1 _21723_ (.A(_12030_),
    .B1(_12033_),
    .B2(_12034_),
    .ZN(_12035_));
 INV_X1 _21724_ (.A(_12023_),
    .ZN(_12036_));
 INV_X1 _21725_ (.A(_12030_),
    .ZN(_12037_));
 OAI211_X1 _21726_ (.A(_12032_),
    .B(_12035_),
    .C1(_12036_),
    .C2(_12037_),
    .ZN(_12038_));
 INV_X1 _21727_ (.A(_12033_),
    .ZN(_12039_));
 INV_X1 _21728_ (.A(_12034_),
    .ZN(_12040_));
 NAND2_X1 _21729_ (.A1(_12039_),
    .A2(_12040_),
    .ZN(_12041_));
 AND2_X1 _21730_ (.A1(_12041_),
    .A2(_12019_),
    .ZN(_12042_));
 NAND2_X1 _21731_ (.A1(_12019_),
    .A2(_11900_),
    .ZN(_12043_));
 INV_X1 _21732_ (.A(_12019_),
    .ZN(_12044_));
 INV_X1 _21733_ (.A(_11894_),
    .ZN(_12045_));
 OAI21_X1 _21734_ (.A(_12043_),
    .B1(_12044_),
    .B2(_12045_),
    .ZN(_12046_));
 NOR4_X1 _21735_ (.A1(_12029_),
    .A2(_12038_),
    .A3(_12042_),
    .A4(_12046_),
    .ZN(_12047_));
 AND2_X1 _21736_ (.A1(_11917_),
    .A2(_11891_),
    .ZN(_12048_));
 NOR2_X2 _21737_ (.A1(_11971_),
    .A2(_16790_),
    .ZN(_12049_));
 AND2_X1 _21738_ (.A1(_12049_),
    .A2(_11924_),
    .ZN(_12050_));
 AND2_X1 _21739_ (.A1(_12048_),
    .A2(_12050_),
    .ZN(_12051_));
 INV_X1 _21740_ (.A(_12051_),
    .ZN(_12052_));
 NAND2_X1 _21741_ (.A1(_11994_),
    .A2(_12050_),
    .ZN(_12053_));
 NAND2_X1 _21742_ (.A1(_11968_),
    .A2(_11904_),
    .ZN(_12054_));
 INV_X1 _21743_ (.A(_12054_),
    .ZN(_12055_));
 NAND2_X1 _21744_ (.A1(_12055_),
    .A2(_12050_),
    .ZN(_12056_));
 AND3_X1 _21745_ (.A1(_12052_),
    .A2(_12053_),
    .A3(_12056_),
    .ZN(_12057_));
 AND2_X1 _21746_ (.A1(_11892_),
    .A2(_11890_),
    .ZN(_12058_));
 AND2_X1 _21747_ (.A1(_12050_),
    .A2(_12058_),
    .ZN(_12059_));
 INV_X1 _21748_ (.A(_12059_),
    .ZN(_12060_));
 OAI211_X1 _21749_ (.A(_12050_),
    .B(_11944_),
    .C1(_11890_),
    .C2(_11933_),
    .ZN(_12061_));
 AND2_X1 _21750_ (.A1(_12060_),
    .A2(_12061_),
    .ZN(_12062_));
 AND2_X1 _21751_ (.A1(_11884_),
    .A2(_12049_),
    .ZN(_12063_));
 BUF_X2 _21752_ (.A(_12063_),
    .Z(_12064_));
 OAI21_X1 _21753_ (.A(_12064_),
    .B1(_12033_),
    .B2(_11955_),
    .ZN(_12065_));
 OAI21_X1 _21754_ (.A(_12064_),
    .B1(_11929_),
    .B2(_11948_),
    .ZN(_12066_));
 AND4_X1 _21755_ (.A1(_12057_),
    .A2(_12062_),
    .A3(_12065_),
    .A4(_12066_),
    .ZN(_12067_));
 AND2_X2 _21756_ (.A1(_11957_),
    .A2(_12049_),
    .ZN(_12068_));
 INV_X2 _21757_ (.A(_12068_),
    .ZN(_12069_));
 INV_X1 _21758_ (.A(_11970_),
    .ZN(_12070_));
 INV_X1 _21759_ (.A(_11980_),
    .ZN(_12071_));
 AOI21_X1 _21760_ (.A(_12069_),
    .B1(_12070_),
    .B2(_12071_),
    .ZN(_12072_));
 NAND2_X1 _21761_ (.A1(_12068_),
    .A2(_11898_),
    .ZN(_12073_));
 NAND3_X1 _21762_ (.A1(_11962_),
    .A2(_11957_),
    .A3(_12049_),
    .ZN(_12074_));
 INV_X1 _21763_ (.A(_12058_),
    .ZN(_12075_));
 OAI211_X1 _21764_ (.A(_12073_),
    .B(_12074_),
    .C1(_12069_),
    .C2(_12075_),
    .ZN(_12076_));
 AND2_X1 _21765_ (.A1(_12049_),
    .A2(_11941_),
    .ZN(_12077_));
 BUF_X2 _21766_ (.A(_12077_),
    .Z(_12078_));
 INV_X2 _21767_ (.A(_12078_),
    .ZN(_12079_));
 AND2_X2 _21768_ (.A1(_11927_),
    .A2(_11893_),
    .ZN(_12080_));
 INV_X1 _21769_ (.A(_12080_),
    .ZN(_12081_));
 AOI21_X1 _21770_ (.A(_12079_),
    .B1(_12081_),
    .B2(_12039_),
    .ZN(_12082_));
 INV_X1 _21771_ (.A(_12001_),
    .ZN(_12083_));
 AND2_X1 _21772_ (.A1(_11904_),
    .A2(_11890_),
    .ZN(_12084_));
 INV_X1 _21773_ (.A(_12084_),
    .ZN(_12085_));
 AOI21_X1 _21774_ (.A(_12079_),
    .B1(_12083_),
    .B2(_12085_),
    .ZN(_12086_));
 NOR4_X1 _21775_ (.A1(_12072_),
    .A2(_12076_),
    .A3(_12082_),
    .A4(_12086_),
    .ZN(_12087_));
 AND2_X2 _21776_ (.A1(_11924_),
    .A2(_12018_),
    .ZN(_12088_));
 BUF_X2 _21777_ (.A(_12088_),
    .Z(_12089_));
 BUF_X2 _21778_ (.A(_12001_),
    .Z(_12090_));
 OAI21_X1 _21779_ (.A(_12089_),
    .B1(_12090_),
    .B2(_11930_),
    .ZN(_12091_));
 AND2_X1 _21780_ (.A1(_11911_),
    .A2(_12018_),
    .ZN(_12092_));
 AND3_X1 _21781_ (.A1(_12092_),
    .A2(_11918_),
    .A3(_11968_),
    .ZN(_12093_));
 BUF_X2 _21782_ (.A(_12092_),
    .Z(_12094_));
 AOI21_X1 _21783_ (.A(_12093_),
    .B1(_12094_),
    .B2(_11953_),
    .ZN(_12095_));
 NOR3_X1 _21784_ (.A1(_11919_),
    .A2(_16786_),
    .A3(_16785_),
    .ZN(_12096_));
 OAI21_X1 _21785_ (.A(_12092_),
    .B1(_11882_),
    .B2(_12096_),
    .ZN(_12097_));
 OAI211_X1 _21786_ (.A(_12089_),
    .B(_11945_),
    .C1(_11955_),
    .C2(_11944_),
    .ZN(_12098_));
 AND4_X1 _21787_ (.A1(_12091_),
    .A2(_12095_),
    .A3(_12097_),
    .A4(_12098_),
    .ZN(_12099_));
 NAND4_X1 _21788_ (.A1(_12047_),
    .A2(_12067_),
    .A3(_12087_),
    .A4(_12099_),
    .ZN(_12100_));
 NOR2_X2 _21789_ (.A1(_12017_),
    .A2(_12100_),
    .ZN(_12101_));
 INV_X2 _21790_ (.A(_12101_),
    .ZN(_12102_));
 XNOR2_X1 _21791_ (.A(_11879_),
    .B(_12102_),
    .ZN(_12103_));
 XNOR2_X1 _21792_ (.A(_12103_),
    .B(_17163_),
    .ZN(_12104_));
 MUX2_X1 _21793_ (.A(_11085_),
    .B(_12104_),
    .S(_11084_),
    .Z(_00716_));
 XOR2_X1 _21794_ (.A(_17174_),
    .B(_16989_),
    .Z(_12105_));
 NAND2_X1 _21795_ (.A1(_11735_),
    .A2(_11604_),
    .ZN(_12106_));
 OAI211_X1 _21796_ (.A(_11750_),
    .B(_12106_),
    .C1(_11739_),
    .C2(_11784_),
    .ZN(_12107_));
 INV_X1 _21797_ (.A(_11674_),
    .ZN(_12108_));
 AOI21_X1 _21798_ (.A(_11739_),
    .B1(_12108_),
    .B2(_11845_),
    .ZN(_12109_));
 AND4_X1 _21799_ (.A1(_11602_),
    .A2(_11709_),
    .A3(_11701_),
    .A4(_11732_),
    .ZN(_12110_));
 NOR3_X1 _21800_ (.A1(_12107_),
    .A2(_12109_),
    .A3(_12110_),
    .ZN(_12111_));
 NAND2_X1 _21801_ (.A1(_11845_),
    .A2(_12108_),
    .ZN(_12112_));
 AND2_X1 _21802_ (.A1(_12112_),
    .A2(_11756_),
    .ZN(_12113_));
 INV_X1 _21803_ (.A(_12113_),
    .ZN(_12114_));
 NAND3_X1 _21804_ (.A1(_11779_),
    .A2(_11732_),
    .A3(_11659_),
    .ZN(_12115_));
 INV_X1 _21805_ (.A(_11756_),
    .ZN(_12116_));
 OAI211_X1 _21806_ (.A(_12114_),
    .B(_12115_),
    .C1(_11811_),
    .C2(_12116_),
    .ZN(_12117_));
 AND2_X1 _21807_ (.A1(_11755_),
    .A2(_11683_),
    .ZN(_12118_));
 AOI21_X1 _21808_ (.A(_11801_),
    .B1(_11684_),
    .B2(_11623_),
    .ZN(_12119_));
 AOI21_X1 _21809_ (.A(_11801_),
    .B1(_11691_),
    .B2(_11840_),
    .ZN(_12120_));
 NOR4_X1 _21810_ (.A1(_12117_),
    .A2(_12118_),
    .A3(_12119_),
    .A4(_12120_),
    .ZN(_12121_));
 BUF_X2 _21811_ (.A(_11743_),
    .Z(_12122_));
 OAI21_X1 _21812_ (.A(_12122_),
    .B1(_11759_),
    .B2(_11598_),
    .ZN(_12123_));
 AND2_X1 _21813_ (.A1(_11674_),
    .A2(_11743_),
    .ZN(_12124_));
 AND2_X1 _21814_ (.A1(_11587_),
    .A2(_12122_),
    .ZN(_12125_));
 AOI211_X1 _21815_ (.A(_12124_),
    .B(_12125_),
    .C1(_11644_),
    .C2(_12122_),
    .ZN(_12126_));
 AND4_X1 _21816_ (.A1(_12111_),
    .A2(_12121_),
    .A3(_12123_),
    .A4(_12126_),
    .ZN(_12127_));
 AOI211_X1 _21817_ (.A(_11568_),
    .B(_11717_),
    .C1(_11707_),
    .C2(_11554_),
    .ZN(_12128_));
 AND2_X1 _21818_ (.A1(_11714_),
    .A2(_11687_),
    .ZN(_12129_));
 AND2_X1 _21819_ (.A1(_11622_),
    .A2(_11713_),
    .ZN(_12130_));
 AND3_X1 _21820_ (.A1(_11713_),
    .A2(_11632_),
    .A3(_11620_),
    .ZN(_12131_));
 NOR4_X1 _21821_ (.A1(_12128_),
    .A2(_12129_),
    .A3(_12130_),
    .A4(_12131_),
    .ZN(_12132_));
 AND2_X1 _21822_ (.A1(_11563_),
    .A2(_11680_),
    .ZN(_12133_));
 AND2_X1 _21823_ (.A1(_11620_),
    .A2(_11824_),
    .ZN(_12134_));
 INV_X1 _21824_ (.A(_12134_),
    .ZN(_12135_));
 OAI21_X1 _21825_ (.A(_11856_),
    .B1(_11692_),
    .B2(_12135_),
    .ZN(_12136_));
 AOI211_X1 _21826_ (.A(_12133_),
    .B(_12136_),
    .C1(_11768_),
    .C2(_11680_),
    .ZN(_12137_));
 OAI21_X1 _21827_ (.A(_11722_),
    .B1(_11720_),
    .B2(_11669_),
    .ZN(_12138_));
 NAND2_X1 _21828_ (.A1(_11598_),
    .A2(_11704_),
    .ZN(_12139_));
 OAI211_X1 _21829_ (.A(_11704_),
    .B(_11571_),
    .C1(_11706_),
    .C2(_11707_),
    .ZN(_12140_));
 OAI211_X1 _21830_ (.A(_11704_),
    .B(_11705_),
    .C1(_11824_),
    .C2(_11559_),
    .ZN(_12141_));
 AND4_X1 _21831_ (.A1(_11700_),
    .A2(_12139_),
    .A3(_12140_),
    .A4(_12141_),
    .ZN(_12142_));
 AND4_X1 _21832_ (.A1(_12132_),
    .A2(_12137_),
    .A3(_12138_),
    .A4(_12142_),
    .ZN(_12143_));
 AOI211_X1 _21833_ (.A(_11786_),
    .B(_11847_),
    .C1(_11671_),
    .C2(_11788_),
    .ZN(_12144_));
 AND2_X1 _21834_ (.A1(_11720_),
    .A2(_11553_),
    .ZN(_12145_));
 AND4_X1 _21835_ (.A1(_11567_),
    .A2(_11566_),
    .A3(_11592_),
    .A4(_11572_),
    .ZN(_12146_));
 AOI21_X1 _21836_ (.A(_11847_),
    .B1(_11811_),
    .B2(_11741_),
    .ZN(_12147_));
 NOR4_X1 _21837_ (.A1(_12144_),
    .A2(_12145_),
    .A3(_12146_),
    .A4(_12147_),
    .ZN(_12148_));
 CLKBUF_X2 _21838_ (.A(_11617_),
    .Z(_12149_));
 NOR2_X1 _21839_ (.A1(_11668_),
    .A2(_11710_),
    .ZN(_12150_));
 AND2_X1 _21840_ (.A1(_12149_),
    .A2(_12150_),
    .ZN(_12151_));
 AOI21_X1 _21841_ (.A(_11618_),
    .B1(_11860_),
    .B2(_11741_),
    .ZN(_12152_));
 AOI211_X1 _21842_ (.A(_12151_),
    .B(_12152_),
    .C1(_12149_),
    .C2(_12134_),
    .ZN(_12153_));
 NAND4_X1 _21843_ (.A1(_11566_),
    .A2(_11672_),
    .A3(_11710_),
    .A4(_11588_),
    .ZN(_12154_));
 OAI21_X1 _21844_ (.A(_12154_),
    .B1(_11591_),
    .B2(_11784_),
    .ZN(_12155_));
 AOI211_X1 _21845_ (.A(_11831_),
    .B(_12155_),
    .C1(_11581_),
    .C2(_11781_),
    .ZN(_12156_));
 AND3_X1 _21846_ (.A1(_11603_),
    .A2(_11788_),
    .A3(_11787_),
    .ZN(_12157_));
 AOI21_X1 _21847_ (.A(_11843_),
    .B1(_11811_),
    .B2(_11780_),
    .ZN(_12158_));
 OR2_X1 _21848_ (.A1(_11833_),
    .A2(_11757_),
    .ZN(_12159_));
 AOI211_X1 _21849_ (.A(_12157_),
    .B(_12158_),
    .C1(_11607_),
    .C2(_12159_),
    .ZN(_12160_));
 AND4_X1 _21850_ (.A1(_12148_),
    .A2(_12153_),
    .A3(_12156_),
    .A4(_12160_),
    .ZN(_12161_));
 AND2_X1 _21851_ (.A1(_11821_),
    .A2(_11749_),
    .ZN(_12162_));
 AND2_X1 _21852_ (.A1(_11664_),
    .A2(_11686_),
    .ZN(_12163_));
 AND2_X1 _21853_ (.A1(_11633_),
    .A2(_11821_),
    .ZN(_12164_));
 AND2_X1 _21854_ (.A1(_11821_),
    .A2(_11627_),
    .ZN(_12165_));
 OR4_X1 _21855_ (.A1(_12162_),
    .A2(_12163_),
    .A3(_12164_),
    .A4(_12165_),
    .ZN(_12166_));
 OAI211_X1 _21856_ (.A(_11656_),
    .B(_11709_),
    .C1(_11701_),
    .C2(_11661_),
    .ZN(_12167_));
 NAND4_X1 _21857_ (.A1(_11701_),
    .A2(_11646_),
    .A3(_11592_),
    .A4(_11572_),
    .ZN(_12168_));
 NAND2_X1 _21858_ (.A1(_11656_),
    .A2(_11609_),
    .ZN(_12169_));
 NAND4_X1 _21859_ (.A1(_12167_),
    .A2(_11651_),
    .A3(_12168_),
    .A4(_12169_),
    .ZN(_12170_));
 AND2_X1 _21860_ (.A1(_11584_),
    .A2(_11582_),
    .ZN(_12171_));
 OAI21_X1 _21861_ (.A(_11675_),
    .B1(_12171_),
    .B2(_11608_),
    .ZN(_12172_));
 AND2_X1 _21862_ (.A1(_11683_),
    .A2(_11667_),
    .ZN(_12173_));
 INV_X1 _21863_ (.A(_12173_),
    .ZN(_12174_));
 OAI211_X1 _21864_ (.A(_12172_),
    .B(_12174_),
    .C1(_11818_),
    .C2(_11654_),
    .ZN(_12175_));
 OAI21_X1 _21865_ (.A(_11639_),
    .B1(_11694_),
    .B2(_11622_),
    .ZN(_12176_));
 NAND2_X1 _21866_ (.A1(_11639_),
    .A2(_11737_),
    .ZN(_12177_));
 OAI211_X1 _21867_ (.A(_12176_),
    .B(_12177_),
    .C1(_11786_),
    .C2(_11783_),
    .ZN(_12178_));
 NOR4_X1 _21868_ (.A1(_12166_),
    .A2(_12170_),
    .A3(_12175_),
    .A4(_12178_),
    .ZN(_12179_));
 NAND4_X1 _21869_ (.A1(_12127_),
    .A2(_12143_),
    .A3(_12161_),
    .A4(_12179_),
    .ZN(_12180_));
 NOR2_X2 _21870_ (.A1(_12180_),
    .A2(_11775_),
    .ZN(_12181_));
 CLKBUF_X2 _21871_ (.A(_11147_),
    .Z(_12182_));
 AND3_X1 _21872_ (.A1(_11215_),
    .A2(_12182_),
    .A3(_11263_),
    .ZN(_12183_));
 AND3_X1 _21873_ (.A1(_11163_),
    .A2(_12182_),
    .A3(_11288_),
    .ZN(_12184_));
 AND2_X1 _21874_ (.A1(_16736_),
    .A2(_16738_),
    .ZN(_12185_));
 NOR2_X1 _21875_ (.A1(_11095_),
    .A2(_16737_),
    .ZN(_12186_));
 AND2_X2 _21876_ (.A1(_12185_),
    .A2(_12186_),
    .ZN(_12187_));
 AOI211_X1 _21877_ (.A(_12183_),
    .B(_12184_),
    .C1(_12187_),
    .C2(_11265_),
    .ZN(_12188_));
 NAND4_X1 _21878_ (.A1(_12182_),
    .A2(_11142_),
    .A3(_11288_),
    .A4(_11239_),
    .ZN(_12189_));
 OAI211_X1 _21879_ (.A(_11265_),
    .B(_11194_),
    .C1(_11150_),
    .C2(_11142_),
    .ZN(_12190_));
 AND3_X1 _21880_ (.A1(_12188_),
    .A2(_12189_),
    .A3(_12190_),
    .ZN(_12191_));
 INV_X1 _21881_ (.A(_11133_),
    .ZN(_12192_));
 AOI21_X1 _21882_ (.A(_11292_),
    .B1(_11280_),
    .B2(_12192_),
    .ZN(_12193_));
 AND2_X1 _21883_ (.A1(_11116_),
    .A2(_11291_),
    .ZN(_12194_));
 AND2_X1 _21884_ (.A1(_11215_),
    .A2(_11291_),
    .ZN(_12195_));
 AND2_X1 _21885_ (.A1(_11217_),
    .A2(_11290_),
    .ZN(_12196_));
 NOR4_X1 _21886_ (.A1(_12193_),
    .A2(_12194_),
    .A3(_12195_),
    .A4(_12196_),
    .ZN(_12197_));
 INV_X1 _21887_ (.A(_11126_),
    .ZN(_12198_));
 NOR2_X1 _21888_ (.A1(_12198_),
    .A2(_11118_),
    .ZN(_12199_));
 AND3_X1 _21889_ (.A1(_11274_),
    .A2(_11203_),
    .A3(_12199_),
    .ZN(_12200_));
 NAND2_X1 _21890_ (.A1(_11274_),
    .A2(_11301_),
    .ZN(_12201_));
 INV_X1 _21891_ (.A(_12187_),
    .ZN(_12202_));
 OAI21_X1 _21892_ (.A(_12201_),
    .B1(_11276_),
    .B2(_12202_),
    .ZN(_12203_));
 AND2_X1 _21893_ (.A1(_11098_),
    .A2(_11118_),
    .ZN(_12204_));
 BUF_X2 _21894_ (.A(_12204_),
    .Z(_12205_));
 AOI211_X1 _21895_ (.A(_12200_),
    .B(_12203_),
    .C1(_12205_),
    .C2(_11285_),
    .ZN(_12206_));
 AND2_X1 _21896_ (.A1(_11282_),
    .A2(_11297_),
    .ZN(_12207_));
 INV_X1 _21897_ (.A(_11297_),
    .ZN(_12208_));
 AOI21_X1 _21898_ (.A(_12208_),
    .B1(_11117_),
    .B2(_11218_),
    .ZN(_12209_));
 AOI211_X1 _21899_ (.A(_12207_),
    .B(_12209_),
    .C1(_12205_),
    .C2(_11299_),
    .ZN(_12210_));
 AND4_X1 _21900_ (.A1(_12191_),
    .A2(_12197_),
    .A3(_12206_),
    .A4(_12210_),
    .ZN(_12211_));
 NAND3_X1 _21901_ (.A1(_11137_),
    .A2(_11184_),
    .A3(_11194_),
    .ZN(_12212_));
 OAI21_X1 _21902_ (.A(_11136_),
    .B1(_11302_),
    .B2(_11304_),
    .ZN(_12213_));
 OAI211_X1 _21903_ (.A(_11136_),
    .B(_11185_),
    .C1(_11125_),
    .C2(_11155_),
    .ZN(_12214_));
 NAND4_X1 _21904_ (.A1(_11091_),
    .A2(_11095_),
    .A3(_11143_),
    .A4(_11153_),
    .ZN(_12215_));
 AND4_X1 _21905_ (.A1(_12212_),
    .A2(_12213_),
    .A3(_12214_),
    .A4(_12215_),
    .ZN(_12216_));
 AND2_X1 _21906_ (.A1(_11092_),
    .A2(_11190_),
    .ZN(_12217_));
 INV_X1 _21907_ (.A(_11092_),
    .ZN(_12218_));
 INV_X1 _21908_ (.A(_11303_),
    .ZN(_12219_));
 AOI21_X1 _21909_ (.A(_12218_),
    .B1(_12219_),
    .B2(_11122_),
    .ZN(_12220_));
 AND2_X1 _21910_ (.A1(_11099_),
    .A2(_11173_),
    .ZN(_12221_));
 AOI211_X1 _21911_ (.A(_12217_),
    .B(_12220_),
    .C1(_11093_),
    .C2(_12221_),
    .ZN(_12222_));
 NAND2_X1 _21912_ (.A1(_11148_),
    .A2(_11301_),
    .ZN(_12223_));
 INV_X1 _21913_ (.A(_11148_),
    .ZN(_12224_));
 OAI21_X1 _21914_ (.A(_12223_),
    .B1(_12224_),
    .B2(_12202_),
    .ZN(_12225_));
 AND2_X1 _21915_ (.A1(_11098_),
    .A2(_11115_),
    .ZN(_12226_));
 INV_X1 _21916_ (.A(_12226_),
    .ZN(_12227_));
 AOI21_X1 _21917_ (.A(_12224_),
    .B1(_11278_),
    .B2(_12227_),
    .ZN(_12228_));
 INV_X1 _21918_ (.A(_11163_),
    .ZN(_12229_));
 NAND2_X1 _21919_ (.A1(_12229_),
    .A2(_11216_),
    .ZN(_12230_));
 AOI211_X1 _21920_ (.A(_12225_),
    .B(_12228_),
    .C1(_11149_),
    .C2(_12230_),
    .ZN(_12231_));
 AND3_X1 _21921_ (.A1(_11225_),
    .A2(_11184_),
    .A3(_11129_),
    .ZN(_12232_));
 NOR2_X1 _21922_ (.A1(_12198_),
    .A2(_11158_),
    .ZN(_12233_));
 AND2_X1 _21923_ (.A1(_12233_),
    .A2(_11103_),
    .ZN(_12234_));
 AND2_X1 _21924_ (.A1(_11103_),
    .A2(_11096_),
    .ZN(_12235_));
 AND4_X1 _21925_ (.A1(_11189_),
    .A2(_11099_),
    .A3(_11091_),
    .A4(_11102_),
    .ZN(_12236_));
 NOR4_X1 _21926_ (.A1(_12232_),
    .A2(_12234_),
    .A3(_12235_),
    .A4(_12236_),
    .ZN(_12237_));
 AND4_X1 _21927_ (.A1(_12216_),
    .A2(_12222_),
    .A3(_12231_),
    .A4(_12237_),
    .ZN(_12238_));
 NOR2_X1 _21928_ (.A1(_11154_),
    .A2(_11125_),
    .ZN(_12239_));
 OAI21_X1 _21929_ (.A(_11221_),
    .B1(_11220_),
    .B2(_12239_),
    .ZN(_12240_));
 AND2_X1 _21930_ (.A1(_11207_),
    .A2(_11160_),
    .ZN(_12241_));
 NAND2_X1 _21931_ (.A1(_11205_),
    .A2(_11303_),
    .ZN(_12242_));
 NAND2_X1 _21932_ (.A1(_11207_),
    .A2(_11121_),
    .ZN(_12243_));
 NAND2_X1 _21933_ (.A1(_12242_),
    .A2(_12243_),
    .ZN(_12244_));
 AOI211_X1 _21934_ (.A(_12241_),
    .B(_12244_),
    .C1(_11207_),
    .C2(_12221_),
    .ZN(_12245_));
 AND2_X1 _21935_ (.A1(_11220_),
    .A2(_11175_),
    .ZN(_12246_));
 AND2_X1 _21936_ (.A1(_11138_),
    .A2(_11171_),
    .ZN(_12247_));
 AND2_X1 _21937_ (.A1(_11175_),
    .A2(_12185_),
    .ZN(_12248_));
 NOR4_X1 _21938_ (.A1(_12246_),
    .A2(_11182_),
    .A3(_12247_),
    .A4(_12248_),
    .ZN(_12249_));
 INV_X1 _21939_ (.A(_11191_),
    .ZN(_12250_));
 INV_X1 _21940_ (.A(_11301_),
    .ZN(_12251_));
 AOI21_X1 _21941_ (.A(_12250_),
    .B1(_12251_),
    .B2(_11117_),
    .ZN(_12252_));
 AOI21_X1 _21942_ (.A(_12250_),
    .B1(_11122_),
    .B2(_11293_),
    .ZN(_12253_));
 AND2_X1 _21943_ (.A1(_11133_),
    .A2(_11191_),
    .ZN(_12254_));
 NOR4_X1 _21944_ (.A1(_12252_),
    .A2(_12253_),
    .A3(_11192_),
    .A4(_12254_),
    .ZN(_12255_));
 AND4_X1 _21945_ (.A1(_12240_),
    .A2(_12245_),
    .A3(_12249_),
    .A4(_12255_),
    .ZN(_12256_));
 INV_X1 _21946_ (.A(_11243_),
    .ZN(_12257_));
 AOI21_X1 _21947_ (.A(_12257_),
    .B1(_11266_),
    .B2(_11122_),
    .ZN(_12258_));
 NAND4_X1 _21948_ (.A1(_11237_),
    .A2(_11173_),
    .A3(_11195_),
    .A4(_11153_),
    .ZN(_12259_));
 INV_X1 _21949_ (.A(_12205_),
    .ZN(_12260_));
 OAI21_X1 _21950_ (.A(_12259_),
    .B1(_12260_),
    .B2(_12257_),
    .ZN(_12261_));
 AND4_X1 _21951_ (.A1(_11095_),
    .A2(_11237_),
    .A3(_11141_),
    .A4(_11195_),
    .ZN(_12262_));
 NOR3_X1 _21952_ (.A1(_12258_),
    .A2(_12261_),
    .A3(_12262_),
    .ZN(_12263_));
 AND2_X1 _21953_ (.A1(_11251_),
    .A2(_11185_),
    .ZN(_12264_));
 NAND2_X1 _21954_ (.A1(_11251_),
    .A2(_11281_),
    .ZN(_12265_));
 INV_X1 _21955_ (.A(_11251_),
    .ZN(_12266_));
 OAI21_X1 _21956_ (.A(_12265_),
    .B1(_12266_),
    .B2(_11268_),
    .ZN(_12267_));
 AOI211_X1 _21957_ (.A(_12264_),
    .B(_12267_),
    .C1(_11302_),
    .C2(_11252_),
    .ZN(_12268_));
 NAND4_X1 _21958_ (.A1(_11231_),
    .A2(_11118_),
    .A3(_11135_),
    .A4(_11153_),
    .ZN(_12269_));
 AND2_X1 _21959_ (.A1(_11233_),
    .A2(_12269_),
    .ZN(_12270_));
 AND2_X1 _21960_ (.A1(_11232_),
    .A2(_11163_),
    .ZN(_12271_));
 INV_X1 _21961_ (.A(_12271_),
    .ZN(_12272_));
 NAND3_X1 _21962_ (.A1(_11234_),
    .A2(_11225_),
    .A3(_11184_),
    .ZN(_12273_));
 AND3_X1 _21963_ (.A1(_12270_),
    .A2(_12272_),
    .A3(_12273_),
    .ZN(_12274_));
 AND2_X2 _21964_ (.A1(_11125_),
    .A2(_11153_),
    .ZN(_12275_));
 NAND2_X1 _21965_ (.A1(_11259_),
    .A2(_12275_),
    .ZN(_12276_));
 AND2_X1 _21966_ (.A1(_11258_),
    .A2(_11166_),
    .ZN(_12277_));
 INV_X1 _21967_ (.A(_12277_),
    .ZN(_12278_));
 NAND2_X1 _21968_ (.A1(_11258_),
    .A2(_11180_),
    .ZN(_12279_));
 NAND2_X1 _21969_ (.A1(_11259_),
    .A2(_11177_),
    .ZN(_12280_));
 AND4_X1 _21970_ (.A1(_12276_),
    .A2(_12278_),
    .A3(_12279_),
    .A4(_12280_),
    .ZN(_12281_));
 AND4_X1 _21971_ (.A1(_12263_),
    .A2(_12268_),
    .A3(_12274_),
    .A4(_12281_),
    .ZN(_12282_));
 NAND4_X1 _21972_ (.A1(_12211_),
    .A2(_12238_),
    .A3(_12256_),
    .A4(_12282_),
    .ZN(_12283_));
 NOR2_X2 _21973_ (.A1(_12283_),
    .A2(_11311_),
    .ZN(_12284_));
 XNOR2_X2 _21974_ (.A(_12181_),
    .B(_12284_),
    .ZN(_12285_));
 XNOR2_X1 _21975_ (.A(_12285_),
    .B(_11878_),
    .ZN(_12286_));
 INV_X1 _21976_ (.A(_11427_),
    .ZN(_12287_));
 INV_X1 _21977_ (.A(_11528_),
    .ZN(_12288_));
 AOI21_X1 _21978_ (.A(_12287_),
    .B1(_11445_),
    .B2(_12288_),
    .ZN(_12289_));
 AND2_X1 _21979_ (.A1(_11410_),
    .A2(_11427_),
    .ZN(_12290_));
 OR4_X1 _21980_ (.A1(_11474_),
    .A2(_12289_),
    .A3(_11428_),
    .A4(_12290_),
    .ZN(_12291_));
 AND2_X1 _21981_ (.A1(_11434_),
    .A2(_11511_),
    .ZN(_12292_));
 OAI21_X1 _21982_ (.A(_11459_),
    .B1(_11410_),
    .B2(_11525_),
    .ZN(_12293_));
 NAND2_X1 _21983_ (.A1(_11436_),
    .A2(_11459_),
    .ZN(_12294_));
 OAI211_X1 _21984_ (.A(_12293_),
    .B(_12294_),
    .C1(_11538_),
    .C2(_11463_),
    .ZN(_12295_));
 AND2_X1 _21985_ (.A1(_11379_),
    .A2(_11333_),
    .ZN(_12296_));
 INV_X1 _21986_ (.A(_12296_),
    .ZN(_12297_));
 NAND2_X1 _21987_ (.A1(_11333_),
    .A2(_11325_),
    .ZN(_12298_));
 AOI21_X1 _21988_ (.A(_11440_),
    .B1(_12297_),
    .B2(_12298_),
    .ZN(_12299_));
 NAND3_X1 _21989_ (.A1(_11370_),
    .A2(_11364_),
    .A3(_11365_),
    .ZN(_12300_));
 NAND3_X1 _21990_ (.A1(_11424_),
    .A2(_11364_),
    .A3(_11365_),
    .ZN(_12301_));
 NAND2_X1 _21991_ (.A1(_12300_),
    .A2(_12301_),
    .ZN(_12302_));
 OR4_X1 _21992_ (.A1(_12292_),
    .A2(_12295_),
    .A3(_12299_),
    .A4(_12302_),
    .ZN(_12303_));
 OAI211_X1 _21993_ (.A(_11415_),
    .B(_11396_),
    .C1(_11338_),
    .C2(_11335_),
    .ZN(_12304_));
 INV_X1 _21994_ (.A(_11530_),
    .ZN(_12305_));
 OAI21_X1 _21995_ (.A(_12304_),
    .B1(_12305_),
    .B2(_11416_),
    .ZN(_12306_));
 NAND3_X1 _21996_ (.A1(_11425_),
    .A2(_11316_),
    .A3(_11365_),
    .ZN(_12307_));
 NAND2_X1 _21997_ (.A1(_11414_),
    .A2(_11473_),
    .ZN(_12308_));
 OAI221_X1 _21998_ (.A(_12307_),
    .B1(_12297_),
    .B2(_11416_),
    .C1(_11472_),
    .C2(_12308_),
    .ZN(_12309_));
 NOR4_X1 _21999_ (.A1(_12291_),
    .A2(_12303_),
    .A3(_12306_),
    .A4(_12309_),
    .ZN(_12310_));
 AND2_X1 _22000_ (.A1(_11488_),
    .A2(_11461_),
    .ZN(_12311_));
 OAI21_X1 _22001_ (.A(_11487_),
    .B1(_11400_),
    .B2(_11398_),
    .ZN(_12312_));
 INV_X1 _22002_ (.A(_11487_),
    .ZN(_12313_));
 OAI21_X1 _22003_ (.A(_12312_),
    .B1(_12313_),
    .B2(_11538_),
    .ZN(_12314_));
 NAND2_X1 _22004_ (.A1(_11340_),
    .A2(_11487_),
    .ZN(_12315_));
 NAND3_X1 _22005_ (.A1(_11487_),
    .A2(_11418_),
    .A3(_11334_),
    .ZN(_12316_));
 NAND2_X1 _22006_ (.A1(_12315_),
    .A2(_12316_),
    .ZN(_12317_));
 INV_X1 _22007_ (.A(_11371_),
    .ZN(_12318_));
 AOI21_X1 _22008_ (.A(_12313_),
    .B1(_12318_),
    .B2(_11526_),
    .ZN(_12319_));
 OR4_X1 _22009_ (.A1(_12311_),
    .A2(_12314_),
    .A3(_12317_),
    .A4(_12319_),
    .ZN(_12320_));
 AND2_X1 _22010_ (.A1(_11333_),
    .A2(_16744_),
    .ZN(_12321_));
 CLKBUF_X2 _22011_ (.A(_12321_),
    .Z(_12322_));
 OAI21_X1 _22012_ (.A(_11536_),
    .B1(_11452_),
    .B2(_12322_),
    .ZN(_12323_));
 AND2_X1 _22013_ (.A1(_11396_),
    .A2(_11360_),
    .ZN(_12324_));
 OAI21_X1 _22014_ (.A(_11536_),
    .B1(_12324_),
    .B2(_11327_),
    .ZN(_12325_));
 NAND2_X1 _22015_ (.A1(_12323_),
    .A2(_12325_),
    .ZN(_12326_));
 OAI21_X1 _22016_ (.A(_11482_),
    .B1(_11511_),
    .B2(_11437_),
    .ZN(_12327_));
 OAI21_X1 _22017_ (.A(_11482_),
    .B1(_11420_),
    .B2(_11321_),
    .ZN(_12328_));
 INV_X1 _22018_ (.A(_11481_),
    .ZN(_12329_));
 OAI211_X1 _22019_ (.A(_12327_),
    .B(_12328_),
    .C1(_12329_),
    .C2(_11443_),
    .ZN(_12330_));
 NAND3_X1 _22020_ (.A1(_11386_),
    .A2(_11335_),
    .A3(_11396_),
    .ZN(_12331_));
 OAI211_X1 _22021_ (.A(_11483_),
    .B(_11373_),
    .C1(_11435_),
    .C2(_11335_),
    .ZN(_12332_));
 OAI211_X1 _22022_ (.A(_11483_),
    .B(_11423_),
    .C1(_11435_),
    .C2(_11472_),
    .ZN(_12333_));
 NAND4_X1 _22023_ (.A1(_11392_),
    .A2(_12331_),
    .A3(_12332_),
    .A4(_12333_),
    .ZN(_12334_));
 NOR4_X1 _22024_ (.A1(_12320_),
    .A2(_12326_),
    .A3(_12330_),
    .A4(_12334_),
    .ZN(_12335_));
 NAND2_X1 _22025_ (.A1(_11542_),
    .A2(_11497_),
    .ZN(_12336_));
 INV_X1 _22026_ (.A(_12298_),
    .ZN(_12337_));
 BUF_X2 _22027_ (.A(_12337_),
    .Z(_12338_));
 OAI21_X1 _22028_ (.A(_11497_),
    .B1(_12338_),
    .B2(_12322_),
    .ZN(_12339_));
 OAI211_X1 _22029_ (.A(_11497_),
    .B(_11423_),
    .C1(_11418_),
    .C2(_11362_),
    .ZN(_12340_));
 NAND4_X1 _22030_ (.A1(_11314_),
    .A2(_11335_),
    .A3(_11389_),
    .A4(_11351_),
    .ZN(_12341_));
 AND4_X1 _22031_ (.A1(_12336_),
    .A2(_12339_),
    .A3(_12340_),
    .A4(_12341_),
    .ZN(_12342_));
 INV_X1 _22032_ (.A(_11390_),
    .ZN(_12343_));
 AND2_X1 _22033_ (.A1(_12343_),
    .A2(_11347_),
    .ZN(_12344_));
 INV_X1 _22034_ (.A(_11331_),
    .ZN(_12345_));
 INV_X1 _22035_ (.A(_11451_),
    .ZN(_12346_));
 INV_X1 _22036_ (.A(_12322_),
    .ZN(_12347_));
 AOI21_X1 _22037_ (.A(_12345_),
    .B1(_12346_),
    .B2(_12347_),
    .ZN(_12348_));
 AOI211_X1 _22038_ (.A(_12344_),
    .B(_12348_),
    .C1(_11347_),
    .C2(_12324_),
    .ZN(_12349_));
 OAI211_X1 _22039_ (.A(_11318_),
    .B(_11373_),
    .C1(_11435_),
    .C2(_11472_),
    .ZN(_12350_));
 OAI21_X1 _22040_ (.A(_11403_),
    .B1(_11467_),
    .B2(_11442_),
    .ZN(_12351_));
 OAI21_X1 _22041_ (.A(_11318_),
    .B1(_11370_),
    .B2(_11425_),
    .ZN(_12352_));
 AND3_X1 _22042_ (.A1(_12350_),
    .A2(_12351_),
    .A3(_12352_),
    .ZN(_12353_));
 AND3_X1 _22043_ (.A1(_11507_),
    .A2(_11408_),
    .A3(_11406_),
    .ZN(_12354_));
 AND2_X1 _22044_ (.A1(_11356_),
    .A2(_11405_),
    .ZN(_12355_));
 AND4_X1 _22045_ (.A1(_11396_),
    .A2(_11314_),
    .A3(_11343_),
    .A4(_11381_),
    .ZN(_12356_));
 NOR4_X1 _22046_ (.A1(_12354_),
    .A2(_12355_),
    .A3(_11531_),
    .A4(_12356_),
    .ZN(_12357_));
 AND4_X1 _22047_ (.A1(_12342_),
    .A2(_12349_),
    .A3(_12353_),
    .A4(_12357_),
    .ZN(_12358_));
 NAND2_X1 _22048_ (.A1(_11380_),
    .A2(_11352_),
    .ZN(_12359_));
 NAND4_X1 _22049_ (.A1(_11368_),
    .A2(_11389_),
    .A3(_11418_),
    .A4(_11351_),
    .ZN(_12360_));
 AND2_X1 _22050_ (.A1(_12359_),
    .A2(_12360_),
    .ZN(_12361_));
 INV_X1 _22051_ (.A(_12361_),
    .ZN(_12362_));
 AND2_X1 _22052_ (.A1(_11353_),
    .A2(_11370_),
    .ZN(_12363_));
 AND3_X1 _22053_ (.A1(_11353_),
    .A2(_11507_),
    .A3(_11408_),
    .ZN(_12364_));
 OR3_X1 _22054_ (.A1(_12362_),
    .A2(_12363_),
    .A3(_12364_),
    .ZN(_12365_));
 BUF_X2 _22055_ (.A(_11477_),
    .Z(_12366_));
 AND2_X1 _22056_ (.A1(_12366_),
    .A2(_11410_),
    .ZN(_12367_));
 AND2_X1 _22057_ (.A1(_11477_),
    .A2(_12337_),
    .ZN(_12368_));
 NOR2_X1 _22058_ (.A1(_12367_),
    .A2(_12368_),
    .ZN(_12369_));
 NAND3_X1 _22059_ (.A1(_11400_),
    .A2(_11364_),
    .A3(_11368_),
    .ZN(_12370_));
 NAND2_X1 _22060_ (.A1(_12366_),
    .A2(_11493_),
    .ZN(_12371_));
 NAND2_X1 _22061_ (.A1(_12366_),
    .A2(_11461_),
    .ZN(_12372_));
 NAND4_X1 _22062_ (.A1(_12369_),
    .A2(_12370_),
    .A3(_12371_),
    .A4(_12372_),
    .ZN(_12373_));
 BUF_X2 _22063_ (.A(_11382_),
    .Z(_12374_));
 BUF_X2 _22064_ (.A(_11429_),
    .Z(_12375_));
 OAI21_X1 _22065_ (.A(_12374_),
    .B1(_12375_),
    .B2(_11452_),
    .ZN(_12376_));
 OAI21_X1 _22066_ (.A(_12374_),
    .B1(_11511_),
    .B2(_11393_),
    .ZN(_12377_));
 NAND4_X1 _22067_ (.A1(_11368_),
    .A2(_11335_),
    .A3(_11373_),
    .A4(_11381_),
    .ZN(_12378_));
 NAND3_X1 _22068_ (.A1(_12376_),
    .A2(_12377_),
    .A3(_12378_),
    .ZN(_12379_));
 OAI21_X1 _22069_ (.A(_11522_),
    .B1(_11420_),
    .B2(_11437_),
    .ZN(_12380_));
 NAND2_X1 _22070_ (.A1(_11522_),
    .A2(_12338_),
    .ZN(_12381_));
 OAI211_X1 _22071_ (.A(_12380_),
    .B(_12381_),
    .C1(_11355_),
    .C2(_11523_),
    .ZN(_12382_));
 NOR4_X1 _22072_ (.A1(_12365_),
    .A2(_12373_),
    .A3(_12379_),
    .A4(_12382_),
    .ZN(_12383_));
 NAND4_X1 _22073_ (.A1(_12310_),
    .A2(_12335_),
    .A3(_12358_),
    .A4(_12383_),
    .ZN(_12384_));
 NOR2_X2 _22074_ (.A1(_12384_),
    .A2(_11449_),
    .ZN(_12385_));
 XNOR2_X1 _22075_ (.A(_12286_),
    .B(_12385_),
    .ZN(_12386_));
 INV_X1 _22076_ (.A(_11964_),
    .ZN(_12387_));
 INV_X1 _22077_ (.A(_12027_),
    .ZN(_12388_));
 NAND2_X1 _22078_ (.A1(_12387_),
    .A2(_12388_),
    .ZN(_12389_));
 AND2_X1 _22079_ (.A1(_12389_),
    .A2(_12022_),
    .ZN(_12390_));
 CLKBUF_X2 _22080_ (.A(_12030_),
    .Z(_12391_));
 NAND3_X1 _22081_ (.A1(_12391_),
    .A2(_11918_),
    .A3(_11927_),
    .ZN(_12392_));
 NAND2_X1 _22082_ (.A1(_12090_),
    .A2(_12391_),
    .ZN(_12393_));
 NOR2_X1 _22083_ (.A1(_12054_),
    .A2(_11909_),
    .ZN(_12394_));
 INV_X1 _22084_ (.A(_12394_),
    .ZN(_12395_));
 OAI211_X1 _22085_ (.A(_12392_),
    .B(_12393_),
    .C1(_12395_),
    .C2(_12037_),
    .ZN(_12396_));
 INV_X1 _22086_ (.A(_11909_),
    .ZN(_12397_));
 NAND2_X1 _22087_ (.A1(_12397_),
    .A2(_11881_),
    .ZN(_12398_));
 NOR2_X1 _22088_ (.A1(_12398_),
    .A2(_11906_),
    .ZN(_12399_));
 INV_X1 _22089_ (.A(_12399_),
    .ZN(_12400_));
 AND2_X2 _22090_ (.A1(_11893_),
    .A2(_16784_),
    .ZN(_12401_));
 INV_X1 _22091_ (.A(_12401_),
    .ZN(_12402_));
 AOI21_X1 _22092_ (.A(_12044_),
    .B1(_12400_),
    .B2(_12402_),
    .ZN(_12403_));
 NAND2_X1 _22093_ (.A1(_12030_),
    .A2(_12401_),
    .ZN(_12404_));
 NAND3_X1 _22094_ (.A1(_12030_),
    .A2(_11927_),
    .A3(_11944_),
    .ZN(_12405_));
 INV_X1 _22095_ (.A(_11882_),
    .ZN(_12406_));
 OAI211_X1 _22096_ (.A(_12404_),
    .B(_12405_),
    .C1(_12406_),
    .C2(_12037_),
    .ZN(_12407_));
 NOR4_X1 _22097_ (.A1(_12390_),
    .A2(_12396_),
    .A3(_12403_),
    .A4(_12407_),
    .ZN(_12408_));
 OAI21_X1 _22098_ (.A(_12094_),
    .B1(_12399_),
    .B2(_12096_),
    .ZN(_12409_));
 CLKBUF_X2 _22099_ (.A(_11907_),
    .Z(_12410_));
 AND2_X1 _22100_ (.A1(_12094_),
    .A2(_12410_),
    .ZN(_12411_));
 BUF_X2 _22101_ (.A(_11948_),
    .Z(_12412_));
 AOI211_X1 _22102_ (.A(_12093_),
    .B(_12411_),
    .C1(_12094_),
    .C2(_12412_),
    .ZN(_12413_));
 BUF_X2 _22103_ (.A(_11944_),
    .Z(_12414_));
 NAND3_X1 _22104_ (.A1(_12089_),
    .A2(_11920_),
    .A3(_12414_),
    .ZN(_12415_));
 NAND2_X1 _22105_ (.A1(_11968_),
    .A2(_11892_),
    .ZN(_12416_));
 INV_X1 _22106_ (.A(_12416_),
    .ZN(_12417_));
 NAND2_X1 _22107_ (.A1(_12417_),
    .A2(_12089_),
    .ZN(_12418_));
 OAI211_X1 _22108_ (.A(_12089_),
    .B(_12011_),
    .C1(_11945_),
    .C2(_11933_),
    .ZN(_12419_));
 NAND2_X1 _22109_ (.A1(_12027_),
    .A2(_12088_),
    .ZN(_12420_));
 AND4_X1 _22110_ (.A1(_12415_),
    .A2(_12418_),
    .A3(_12419_),
    .A4(_12420_),
    .ZN(_12421_));
 AND4_X1 _22111_ (.A1(_12408_),
    .A2(_12409_),
    .A3(_12413_),
    .A4(_12421_),
    .ZN(_12422_));
 BUF_X2 _22112_ (.A(_12063_),
    .Z(_12423_));
 OAI21_X1 _22113_ (.A(_12423_),
    .B1(_12058_),
    .B2(_12414_),
    .ZN(_12424_));
 AND2_X1 _22114_ (.A1(_11918_),
    .A2(_11890_),
    .ZN(_12425_));
 INV_X1 _22115_ (.A(_12425_),
    .ZN(_12426_));
 AOI21_X1 _22116_ (.A(_12069_),
    .B1(_12071_),
    .B2(_12426_),
    .ZN(_12427_));
 NAND2_X1 _22117_ (.A1(_12068_),
    .A2(_11882_),
    .ZN(_12428_));
 INV_X1 _22118_ (.A(_11891_),
    .ZN(_12429_));
 NAND2_X1 _22119_ (.A1(_12429_),
    .A2(_11893_),
    .ZN(_12430_));
 OAI21_X1 _22120_ (.A(_12428_),
    .B1(_12069_),
    .B2(_12430_),
    .ZN(_12431_));
 INV_X1 _22121_ (.A(_11900_),
    .ZN(_12432_));
 AOI21_X1 _22122_ (.A(_12079_),
    .B1(_12432_),
    .B2(_12040_),
    .ZN(_12433_));
 OAI21_X1 _22123_ (.A(_12078_),
    .B1(_12003_),
    .B2(_12024_),
    .ZN(_12434_));
 NAND4_X1 _22124_ (.A1(_11918_),
    .A2(_12049_),
    .A3(_11890_),
    .A4(_11941_),
    .ZN(_12435_));
 NAND2_X1 _22125_ (.A1(_12434_),
    .A2(_12435_),
    .ZN(_12436_));
 NOR4_X1 _22126_ (.A1(_12427_),
    .A2(_12431_),
    .A3(_12433_),
    .A4(_12436_),
    .ZN(_12437_));
 NOR3_X1 _22127_ (.A1(_11920_),
    .A2(_11916_),
    .A3(_16785_),
    .ZN(_12438_));
 OAI21_X1 _22128_ (.A(_12423_),
    .B1(_12438_),
    .B2(_12003_),
    .ZN(_12439_));
 BUF_X2 _22129_ (.A(_12050_),
    .Z(_12440_));
 NAND3_X1 _22130_ (.A1(_12055_),
    .A2(_12397_),
    .A3(_12440_),
    .ZN(_12441_));
 NAND2_X1 _22131_ (.A1(_11964_),
    .A2(_12440_),
    .ZN(_12442_));
 NAND2_X1 _22132_ (.A1(_12441_),
    .A2(_12442_),
    .ZN(_12443_));
 NAND2_X1 _22133_ (.A1(_12080_),
    .A2(_12440_),
    .ZN(_12444_));
 INV_X1 _22134_ (.A(_12050_),
    .ZN(_12445_));
 OAI21_X1 _22135_ (.A(_12444_),
    .B1(_12445_),
    .B2(_11988_),
    .ZN(_12446_));
 BUF_X2 _22136_ (.A(_11985_),
    .Z(_12447_));
 AND2_X1 _22137_ (.A1(_12440_),
    .A2(_12447_),
    .ZN(_12448_));
 AND2_X1 _22138_ (.A1(_11881_),
    .A2(_11890_),
    .ZN(_12449_));
 AND2_X1 _22139_ (.A1(_12449_),
    .A2(_12440_),
    .ZN(_12450_));
 NOR4_X1 _22140_ (.A1(_12443_),
    .A2(_12446_),
    .A3(_12448_),
    .A4(_12450_),
    .ZN(_12451_));
 AND4_X1 _22141_ (.A1(_12424_),
    .A2(_12437_),
    .A3(_12439_),
    .A4(_12451_),
    .ZN(_12452_));
 AND2_X1 _22142_ (.A1(_12014_),
    .A2(_11983_),
    .ZN(_12453_));
 AOI21_X1 _22143_ (.A(_11984_),
    .B1(_12054_),
    .B2(_12426_),
    .ZN(_12454_));
 AND2_X1 _22144_ (.A1(_11893_),
    .A2(_11896_),
    .ZN(_12455_));
 AOI211_X1 _22145_ (.A(_12453_),
    .B(_12454_),
    .C1(_11993_),
    .C2(_12455_),
    .ZN(_12456_));
 AND2_X1 _22146_ (.A1(_12000_),
    .A2(_11907_),
    .ZN(_12457_));
 INV_X1 _22147_ (.A(_12000_),
    .ZN(_12458_));
 NOR2_X1 _22148_ (.A1(_12401_),
    .A2(_12455_),
    .ZN(_12459_));
 NOR2_X1 _22149_ (.A1(_12458_),
    .A2(_12459_),
    .ZN(_12460_));
 BUF_X2 _22150_ (.A(_12000_),
    .Z(_12461_));
 AOI211_X1 _22151_ (.A(_12457_),
    .B(_12460_),
    .C1(_12461_),
    .C2(_12014_),
    .ZN(_12462_));
 AND3_X1 _22152_ (.A1(_11974_),
    .A2(_12417_),
    .A3(_12397_),
    .ZN(_12463_));
 AOI21_X1 _22153_ (.A(_12463_),
    .B1(_12412_),
    .B2(_11974_),
    .ZN(_12464_));
 OAI211_X1 _22154_ (.A(_11911_),
    .B(_11979_),
    .C1(_11980_),
    .C2(_12024_),
    .ZN(_12465_));
 NAND3_X1 _22155_ (.A1(_11929_),
    .A2(_11911_),
    .A3(_11979_),
    .ZN(_12466_));
 NAND2_X1 _22156_ (.A1(_12006_),
    .A2(_12034_),
    .ZN(_12467_));
 AND3_X1 _22157_ (.A1(_12465_),
    .A2(_12466_),
    .A3(_12467_),
    .ZN(_12468_));
 AND4_X1 _22158_ (.A1(_12456_),
    .A2(_12462_),
    .A3(_12464_),
    .A4(_12468_),
    .ZN(_12469_));
 AND2_X1 _22159_ (.A1(_11894_),
    .A2(_11943_),
    .ZN(_12470_));
 AND2_X1 _22160_ (.A1(_12425_),
    .A2(_11943_),
    .ZN(_12471_));
 AND3_X1 _22161_ (.A1(_11942_),
    .A2(_11920_),
    .A3(_12011_),
    .ZN(_12472_));
 AND2_X1 _22162_ (.A1(_12024_),
    .A2(_11942_),
    .ZN(_12473_));
 NOR4_X1 _22163_ (.A1(_12470_),
    .A2(_12471_),
    .A3(_12472_),
    .A4(_12473_),
    .ZN(_12474_));
 INV_X1 _22164_ (.A(_11887_),
    .ZN(_12475_));
 NOR3_X1 _22165_ (.A1(_12475_),
    .A2(_11927_),
    .A3(_12430_),
    .ZN(_12476_));
 AND2_X1 _22166_ (.A1(_11887_),
    .A2(_12084_),
    .ZN(_12477_));
 AND2_X1 _22167_ (.A1(_11887_),
    .A2(_11937_),
    .ZN(_12478_));
 NOR4_X1 _22168_ (.A1(_11923_),
    .A2(_12476_),
    .A3(_12477_),
    .A4(_12478_),
    .ZN(_12479_));
 BUF_X2 _22169_ (.A(_11959_),
    .Z(_12480_));
 INV_X1 _22170_ (.A(_12480_),
    .ZN(_12481_));
 OAI21_X1 _22171_ (.A(_11960_),
    .B1(_12481_),
    .B2(_11991_),
    .ZN(_12482_));
 AND3_X1 _22172_ (.A1(_12055_),
    .A2(_11959_),
    .A3(_12397_),
    .ZN(_12483_));
 AND2_X1 _22173_ (.A1(_12480_),
    .A2(_12090_),
    .ZN(_12484_));
 AND2_X1 _22174_ (.A1(_11959_),
    .A2(_11994_),
    .ZN(_12485_));
 NOR4_X1 _22175_ (.A1(_12482_),
    .A2(_12483_),
    .A3(_12484_),
    .A4(_12485_),
    .ZN(_12486_));
 AND2_X1 _22176_ (.A1(_12034_),
    .A2(_11926_),
    .ZN(_12487_));
 INV_X1 _22177_ (.A(_12487_),
    .ZN(_12488_));
 BUF_X2 _22178_ (.A(_11926_),
    .Z(_12489_));
 NAND2_X1 _22179_ (.A1(_12003_),
    .A2(_12489_),
    .ZN(_12490_));
 OAI211_X1 _22180_ (.A(_11926_),
    .B(_11955_),
    .C1(_11945_),
    .C2(_11946_),
    .ZN(_12491_));
 OAI21_X1 _22181_ (.A(_11926_),
    .B1(_12090_),
    .B2(_11994_),
    .ZN(_12492_));
 AND4_X1 _22182_ (.A1(_12488_),
    .A2(_12490_),
    .A3(_12491_),
    .A4(_12492_),
    .ZN(_12493_));
 AND4_X1 _22183_ (.A1(_12474_),
    .A2(_12479_),
    .A3(_12486_),
    .A4(_12493_),
    .ZN(_12494_));
 NAND4_X1 _22184_ (.A1(_12422_),
    .A2(_12452_),
    .A3(_12469_),
    .A4(_12494_),
    .ZN(_12495_));
 OAI21_X1 _22185_ (.A(_11916_),
    .B1(_11968_),
    .B2(_16785_),
    .ZN(_12496_));
 AND3_X1 _22186_ (.A1(_12018_),
    .A2(_11941_),
    .A3(_11916_),
    .ZN(_12497_));
 AND2_X1 _22187_ (.A1(_12496_),
    .A2(_12497_),
    .ZN(_12498_));
 NOR2_X2 _22188_ (.A1(_12495_),
    .A2(_12498_),
    .ZN(_12499_));
 XNOR2_X2 _22189_ (.A(_12499_),
    .B(_12102_),
    .ZN(_12500_));
 XNOR2_X1 _22190_ (.A(_12386_),
    .B(_12500_),
    .ZN(_12501_));
 XNOR2_X1 _22191_ (.A(_12501_),
    .B(_17174_),
    .ZN(_12502_));
 MUX2_X1 _22192_ (.A(_12105_),
    .B(_12502_),
    .S(_11084_),
    .Z(_00717_));
 XOR2_X1 _22193_ (.A(_17185_),
    .B(_16990_),
    .Z(_12503_));
 NOR2_X1 _22194_ (.A1(_11563_),
    .A2(_11587_),
    .ZN(_12504_));
 INV_X1 _22195_ (.A(_12504_),
    .ZN(_12505_));
 BUF_X2 _22196_ (.A(_11867_),
    .Z(_12506_));
 NOR2_X1 _22197_ (.A1(_11689_),
    .A2(_12506_),
    .ZN(_12507_));
 INV_X1 _22198_ (.A(_12507_),
    .ZN(_12508_));
 OAI21_X1 _22199_ (.A(_12149_),
    .B1(_12505_),
    .B2(_12508_),
    .ZN(_12509_));
 AND2_X1 _22200_ (.A1(_12149_),
    .A2(_11627_),
    .ZN(_12510_));
 AND2_X1 _22201_ (.A1(_12149_),
    .A2(_11749_),
    .ZN(_12511_));
 AOI211_X1 _22202_ (.A(_12510_),
    .B(_12511_),
    .C1(_11833_),
    .C2(_12149_),
    .ZN(_12512_));
 OAI21_X1 _22203_ (.A(_11581_),
    .B1(_12506_),
    .B2(_11737_),
    .ZN(_12513_));
 OAI21_X1 _22204_ (.A(_11581_),
    .B1(_11598_),
    .B2(_11612_),
    .ZN(_12514_));
 AND4_X1 _22205_ (.A1(_12509_),
    .A2(_12512_),
    .A3(_12513_),
    .A4(_12514_),
    .ZN(_12515_));
 OAI21_X1 _22206_ (.A(_11553_),
    .B1(_11749_),
    .B2(_11694_),
    .ZN(_12516_));
 OAI21_X1 _22207_ (.A(_11553_),
    .B1(_11779_),
    .B2(_11644_),
    .ZN(_12517_));
 OAI21_X1 _22208_ (.A(_11607_),
    .B1(_11749_),
    .B2(_11612_),
    .ZN(_12518_));
 OAI21_X1 _22209_ (.A(_11607_),
    .B1(_11779_),
    .B2(_11762_),
    .ZN(_12519_));
 AND4_X1 _22210_ (.A1(_12516_),
    .A2(_12517_),
    .A3(_12518_),
    .A4(_12519_),
    .ZN(_12520_));
 AOI21_X1 _22211_ (.A(_11564_),
    .B1(_11709_),
    .B2(_11671_),
    .ZN(_12521_));
 NOR2_X1 _22212_ (.A1(_11683_),
    .A2(_11612_),
    .ZN(_12522_));
 AOI21_X1 _22213_ (.A(_11692_),
    .B1(_12521_),
    .B2(_12522_),
    .ZN(_12523_));
 OAI21_X1 _22214_ (.A(_11714_),
    .B1(_11609_),
    .B2(_11564_),
    .ZN(_12524_));
 OAI21_X1 _22215_ (.A(_12524_),
    .B1(_11780_),
    .B2(_11717_),
    .ZN(_12525_));
 AND2_X1 _22216_ (.A1(_11604_),
    .A2(_11714_),
    .ZN(_12526_));
 AND3_X1 _22217_ (.A1(_11640_),
    .A2(_11582_),
    .A3(_11714_),
    .ZN(_12527_));
 NOR4_X1 _22218_ (.A1(_12523_),
    .A2(_12525_),
    .A3(_12526_),
    .A4(_12527_),
    .ZN(_12528_));
 NOR2_X1 _22219_ (.A1(_11668_),
    .A2(_11701_),
    .ZN(_12529_));
 NAND2_X1 _22220_ (.A1(_11722_),
    .A2(_12529_),
    .ZN(_12530_));
 INV_X1 _22221_ (.A(_11721_),
    .ZN(_12531_));
 OAI211_X1 _22222_ (.A(_11866_),
    .B(_12530_),
    .C1(_11623_),
    .C2(_12531_),
    .ZN(_12532_));
 INV_X1 _22223_ (.A(_11685_),
    .ZN(_12533_));
 AOI21_X1 _22224_ (.A(_11872_),
    .B1(_12533_),
    .B2(_11595_),
    .ZN(_12534_));
 INV_X1 _22225_ (.A(_11689_),
    .ZN(_12535_));
 AOI21_X1 _22226_ (.A(_11872_),
    .B1(_12535_),
    .B2(_11850_),
    .ZN(_12536_));
 NAND2_X1 _22227_ (.A1(_11722_),
    .A2(_11737_),
    .ZN(_12537_));
 NAND3_X1 _22228_ (.A1(_11779_),
    .A2(_11695_),
    .A3(_11659_),
    .ZN(_12538_));
 OAI211_X1 _22229_ (.A(_12537_),
    .B(_12538_),
    .C1(_12531_),
    .C2(_11845_),
    .ZN(_12539_));
 NOR4_X1 _22230_ (.A1(_12532_),
    .A2(_12534_),
    .A3(_12536_),
    .A4(_12539_),
    .ZN(_12540_));
 NAND4_X1 _22231_ (.A1(_12515_),
    .A2(_12520_),
    .A3(_12528_),
    .A4(_12540_),
    .ZN(_12541_));
 OAI21_X1 _22232_ (.A(_11821_),
    .B1(_12171_),
    .B2(_11779_),
    .ZN(_12542_));
 NAND2_X1 _22233_ (.A1(_11821_),
    .A2(_11749_),
    .ZN(_12543_));
 INV_X1 _22234_ (.A(_11664_),
    .ZN(_12544_));
 OAI211_X1 _22235_ (.A(_12542_),
    .B(_12543_),
    .C1(_11619_),
    .C2(_12544_),
    .ZN(_12545_));
 AND2_X1 _22236_ (.A1(_11622_),
    .A2(_11675_),
    .ZN(_12546_));
 OR3_X1 _22237_ (.A1(_12546_),
    .A2(_12173_),
    .A3(_11670_),
    .ZN(_12547_));
 AOI21_X1 _22238_ (.A(_11818_),
    .B1(_11780_),
    .B2(_11811_),
    .ZN(_12548_));
 AND4_X1 _22239_ (.A1(_11824_),
    .A2(_11646_),
    .A3(_11705_),
    .A4(_11588_),
    .ZN(_12549_));
 NOR4_X1 _22240_ (.A1(_12545_),
    .A2(_12547_),
    .A3(_12548_),
    .A4(_12549_),
    .ZN(_12550_));
 OAI21_X1 _22241_ (.A(_11656_),
    .B1(_11604_),
    .B2(_11622_),
    .ZN(_12551_));
 NOR2_X1 _22242_ (.A1(_12521_),
    .A2(_11783_),
    .ZN(_12552_));
 AOI21_X1 _22243_ (.A(_12552_),
    .B1(_11639_),
    .B2(_11687_),
    .ZN(_12553_));
 OAI21_X1 _22244_ (.A(_11650_),
    .B1(_11612_),
    .B2(_11577_),
    .ZN(_12554_));
 OAI211_X1 _22245_ (.A(_11656_),
    .B(_16698_),
    .C1(_11707_),
    .C2(_11554_),
    .ZN(_12555_));
 AND4_X1 _22246_ (.A1(_12551_),
    .A2(_12553_),
    .A3(_12554_),
    .A4(_12555_),
    .ZN(_12556_));
 OAI21_X1 _22247_ (.A(_11756_),
    .B1(_11781_),
    .B2(_11787_),
    .ZN(_12557_));
 OAI21_X1 _22248_ (.A(_11767_),
    .B1(_11768_),
    .B2(_11762_),
    .ZN(_12558_));
 OAI21_X1 _22249_ (.A(_11767_),
    .B1(_11759_),
    .B2(_11622_),
    .ZN(_12559_));
 AND4_X1 _22250_ (.A1(_11804_),
    .A2(_12557_),
    .A3(_12558_),
    .A4(_12559_),
    .ZN(_12560_));
 OAI211_X1 _22251_ (.A(_12122_),
    .B(_11709_),
    .C1(_11706_),
    .C2(_11642_),
    .ZN(_12561_));
 NAND2_X1 _22252_ (.A1(_12506_),
    .A2(_12122_),
    .ZN(_12562_));
 NAND2_X1 _22253_ (.A1(_12561_),
    .A2(_12562_),
    .ZN(_12563_));
 INV_X1 _22254_ (.A(_12563_),
    .ZN(_12564_));
 OAI211_X1 _22255_ (.A(_11735_),
    .B(_11709_),
    .C1(_11701_),
    .C2(_11661_),
    .ZN(_12565_));
 NAND3_X1 _22256_ (.A1(_11674_),
    .A2(_11602_),
    .A3(_11732_),
    .ZN(_12566_));
 NAND2_X1 _22257_ (.A1(_11734_),
    .A2(_11643_),
    .ZN(_12567_));
 AND3_X1 _22258_ (.A1(_12565_),
    .A2(_12566_),
    .A3(_12567_),
    .ZN(_12568_));
 OAI21_X1 _22259_ (.A(_12122_),
    .B1(_11687_),
    .B2(_11702_),
    .ZN(_12569_));
 NAND2_X1 _22260_ (.A1(_11627_),
    .A2(_11735_),
    .ZN(_12570_));
 NAND2_X1 _22261_ (.A1(_11735_),
    .A2(_11687_),
    .ZN(_12571_));
 AND3_X1 _22262_ (.A1(_12106_),
    .A2(_12570_),
    .A3(_12571_),
    .ZN(_12572_));
 AND4_X1 _22263_ (.A1(_12564_),
    .A2(_12568_),
    .A3(_12569_),
    .A4(_12572_),
    .ZN(_12573_));
 NAND4_X1 _22264_ (.A1(_12550_),
    .A2(_12556_),
    .A3(_12560_),
    .A4(_12573_),
    .ZN(_12574_));
 NOR2_X2 _22265_ (.A1(_12541_),
    .A2(_12574_),
    .ZN(_12575_));
 AND2_X1 _22266_ (.A1(_11152_),
    .A2(_11265_),
    .ZN(_12576_));
 AND2_X1 _22267_ (.A1(_12275_),
    .A2(_11265_),
    .ZN(_12577_));
 AOI211_X1 _22268_ (.A(_12576_),
    .B(_12577_),
    .C1(_11181_),
    .C2(_11265_),
    .ZN(_12578_));
 AND2_X1 _22269_ (.A1(_11264_),
    .A2(_11235_),
    .ZN(_12579_));
 AND2_X1 _22270_ (.A1(_11225_),
    .A2(_11183_),
    .ZN(_12580_));
 AOI211_X1 _22271_ (.A(_12183_),
    .B(_12579_),
    .C1(_11265_),
    .C2(_12580_),
    .ZN(_12581_));
 OAI21_X1 _22272_ (.A(_11295_),
    .B1(_11181_),
    .B2(_11100_),
    .ZN(_12582_));
 OAI211_X1 _22273_ (.A(_11295_),
    .B(_11141_),
    .C1(_11150_),
    .C2(_11142_),
    .ZN(_12583_));
 NAND2_X1 _22274_ (.A1(_11128_),
    .A2(_11295_),
    .ZN(_12584_));
 NAND2_X1 _22275_ (.A1(_12583_),
    .A2(_12584_),
    .ZN(_12585_));
 INV_X1 _22276_ (.A(_12585_),
    .ZN(_12586_));
 AND4_X1 _22277_ (.A1(_12578_),
    .A2(_12581_),
    .A3(_12582_),
    .A4(_12586_),
    .ZN(_12587_));
 INV_X1 _22278_ (.A(_11259_),
    .ZN(_12588_));
 INV_X1 _22279_ (.A(_11151_),
    .ZN(_12589_));
 OAI21_X1 _22280_ (.A(_12280_),
    .B1(_12588_),
    .B2(_12589_),
    .ZN(_12590_));
 AND2_X1 _22281_ (.A1(_11259_),
    .A2(_12187_),
    .ZN(_12591_));
 AND3_X1 _22282_ (.A1(_11259_),
    .A2(_12233_),
    .A3(_11184_),
    .ZN(_12592_));
 NOR3_X1 _22283_ (.A1(_12590_),
    .A2(_12591_),
    .A3(_12592_),
    .ZN(_12593_));
 OAI21_X1 _22284_ (.A(_11247_),
    .B1(_12205_),
    .B2(_11282_),
    .ZN(_12594_));
 OAI21_X1 _22285_ (.A(_11247_),
    .B1(_11302_),
    .B2(_12187_),
    .ZN(_12595_));
 NAND4_X1 _22286_ (.A1(_11238_),
    .A2(_11185_),
    .A3(_11195_),
    .A4(_11173_),
    .ZN(_12596_));
 AND2_X1 _22287_ (.A1(_12595_),
    .A2(_12596_),
    .ZN(_12597_));
 AND4_X1 _22288_ (.A1(_11249_),
    .A2(_12593_),
    .A3(_12594_),
    .A4(_12597_),
    .ZN(_12598_));
 OAI21_X1 _22289_ (.A(_11299_),
    .B1(_11304_),
    .B2(_11286_),
    .ZN(_12599_));
 OAI21_X1 _22290_ (.A(_11285_),
    .B1(_12580_),
    .B2(_12199_),
    .ZN(_12600_));
 OAI21_X1 _22291_ (.A(_11299_),
    .B1(_11279_),
    .B2(_11282_),
    .ZN(_12601_));
 NAND3_X1 _22292_ (.A1(_11152_),
    .A2(_11255_),
    .A3(_11288_),
    .ZN(_12602_));
 AND4_X1 _22293_ (.A1(_12599_),
    .A2(_12600_),
    .A3(_12601_),
    .A4(_12602_),
    .ZN(_12603_));
 OAI21_X1 _22294_ (.A(_11252_),
    .B1(_11302_),
    .B2(_11116_),
    .ZN(_12604_));
 NAND2_X1 _22295_ (.A1(_11251_),
    .A2(_11180_),
    .ZN(_12605_));
 OAI211_X1 _22296_ (.A(_12604_),
    .B(_12605_),
    .C1(_11293_),
    .C2(_12266_),
    .ZN(_12606_));
 INV_X1 _22297_ (.A(_11232_),
    .ZN(_12607_));
 AOI21_X1 _22298_ (.A(_12607_),
    .B1(_11277_),
    .B2(_11111_),
    .ZN(_12608_));
 NAND2_X1 _22299_ (.A1(_11234_),
    .A2(_11302_),
    .ZN(_12609_));
 NAND2_X1 _22300_ (.A1(_11234_),
    .A2(_11304_),
    .ZN(_12610_));
 NAND3_X1 _22301_ (.A1(_11139_),
    .A2(_11238_),
    .A3(_11143_),
    .ZN(_12611_));
 NAND3_X1 _22302_ (.A1(_12609_),
    .A2(_12610_),
    .A3(_12611_),
    .ZN(_12612_));
 AND3_X1 _22303_ (.A1(_11238_),
    .A2(_11100_),
    .A3(_11143_),
    .ZN(_12613_));
 NOR4_X1 _22304_ (.A1(_12606_),
    .A2(_12608_),
    .A3(_12612_),
    .A4(_12613_),
    .ZN(_12614_));
 NAND4_X1 _22305_ (.A1(_12587_),
    .A2(_12598_),
    .A3(_12603_),
    .A4(_12614_),
    .ZN(_12615_));
 INV_X1 _22306_ (.A(_11204_),
    .ZN(_12616_));
 AND2_X1 _22307_ (.A1(_12233_),
    .A2(_11183_),
    .ZN(_12617_));
 INV_X1 _22308_ (.A(_12617_),
    .ZN(_12618_));
 AOI21_X1 _22309_ (.A(_12218_),
    .B1(_12616_),
    .B2(_12618_),
    .ZN(_12619_));
 NAND2_X1 _22310_ (.A1(_11129_),
    .A2(_11133_),
    .ZN(_12620_));
 NAND2_X1 _22311_ (.A1(_12620_),
    .A2(_11106_),
    .ZN(_12621_));
 AOI21_X1 _22312_ (.A(_11107_),
    .B1(_11266_),
    .B2(_12251_),
    .ZN(_12622_));
 INV_X1 _22313_ (.A(_12275_),
    .ZN(_12623_));
 AOI21_X1 _22314_ (.A(_12218_),
    .B1(_12623_),
    .B2(_12192_),
    .ZN(_12624_));
 NOR4_X1 _22315_ (.A1(_12619_),
    .A2(_12621_),
    .A3(_12622_),
    .A4(_12624_),
    .ZN(_12625_));
 OAI21_X1 _22316_ (.A(_11137_),
    .B1(_11177_),
    .B2(_11267_),
    .ZN(_12626_));
 OAI21_X1 _22317_ (.A(_11149_),
    .B1(_11177_),
    .B2(_11105_),
    .ZN(_12627_));
 OAI21_X1 _22318_ (.A(_11137_),
    .B1(_12187_),
    .B2(_11235_),
    .ZN(_12628_));
 OAI21_X1 _22319_ (.A(_11149_),
    .B1(_12187_),
    .B2(_11286_),
    .ZN(_12629_));
 AND4_X1 _22320_ (.A1(_12626_),
    .A2(_12627_),
    .A3(_12628_),
    .A4(_12629_),
    .ZN(_12630_));
 AOI22_X1 _22321_ (.A1(_11270_),
    .A2(_11185_),
    .B1(_12186_),
    .B2(_12185_),
    .ZN(_12631_));
 NAND2_X1 _22322_ (.A1(_11190_),
    .A2(_11175_),
    .ZN(_12632_));
 OAI221_X1 _22323_ (.A(_11176_),
    .B1(_12631_),
    .B2(_11172_),
    .C1(_11115_),
    .C2(_12632_),
    .ZN(_12633_));
 AOI21_X1 _22324_ (.A(_11209_),
    .B1(_11277_),
    .B2(_12260_),
    .ZN(_12634_));
 AND3_X1 _22325_ (.A1(_11139_),
    .A2(_11193_),
    .A3(_12182_),
    .ZN(_12635_));
 AOI21_X1 _22326_ (.A(_11209_),
    .B1(_12251_),
    .B2(_11117_),
    .ZN(_12636_));
 NOR4_X1 _22327_ (.A1(_12633_),
    .A2(_12634_),
    .A3(_12635_),
    .A4(_12636_),
    .ZN(_12637_));
 AOI21_X1 _22328_ (.A(_11214_),
    .B1(_12589_),
    .B2(_11283_),
    .ZN(_12638_));
 NAND4_X1 _22329_ (.A1(_11255_),
    .A2(_11193_),
    .A3(_12185_),
    .A4(_12186_),
    .ZN(_12639_));
 NAND4_X1 _22330_ (.A1(_11255_),
    .A2(_11115_),
    .A3(_11185_),
    .A4(_11193_),
    .ZN(_12640_));
 OAI211_X1 _22331_ (.A(_12639_),
    .B(_12640_),
    .C1(_11214_),
    .C2(_12251_),
    .ZN(_12641_));
 AND2_X1 _22332_ (.A1(_11141_),
    .A2(_11189_),
    .ZN(_12642_));
 OAI21_X1 _22333_ (.A(_11199_),
    .B1(_12642_),
    .B2(_11286_),
    .ZN(_12643_));
 NAND4_X1 _22334_ (.A1(_11195_),
    .A2(_11193_),
    .A3(_11239_),
    .A4(_11109_),
    .ZN(_12644_));
 NAND4_X1 _22335_ (.A1(_11199_),
    .A2(_11184_),
    .A3(_11186_),
    .A4(_11100_),
    .ZN(_12645_));
 NAND3_X1 _22336_ (.A1(_12643_),
    .A2(_12644_),
    .A3(_12645_),
    .ZN(_12646_));
 AND2_X1 _22337_ (.A1(_11221_),
    .A2(_11156_),
    .ZN(_12647_));
 NOR4_X1 _22338_ (.A1(_12638_),
    .A2(_12641_),
    .A3(_12646_),
    .A4(_12647_),
    .ZN(_12648_));
 NAND4_X1 _22339_ (.A1(_12625_),
    .A2(_12630_),
    .A3(_12637_),
    .A4(_12648_),
    .ZN(_12649_));
 NOR2_X2 _22340_ (.A1(_12615_),
    .A2(_12649_),
    .ZN(_12650_));
 XOR2_X2 _22341_ (.A(_12575_),
    .B(_12650_),
    .Z(_12651_));
 AND2_X1 _22342_ (.A1(_11382_),
    .A2(_11451_),
    .ZN(_12652_));
 NAND2_X1 _22343_ (.A1(_11521_),
    .A2(_11461_),
    .ZN(_12653_));
 NAND2_X1 _22344_ (.A1(_12653_),
    .A2(_12381_),
    .ZN(_12654_));
 AOI211_X1 _22345_ (.A(_12652_),
    .B(_12654_),
    .C1(_12296_),
    .C2(_11403_),
    .ZN(_12655_));
 AND2_X1 _22346_ (.A1(_11518_),
    .A2(_11488_),
    .ZN(_12656_));
 AND3_X1 _22347_ (.A1(_11534_),
    .A2(_11376_),
    .A3(_11319_),
    .ZN(_12657_));
 AND2_X1 _22348_ (.A1(_12322_),
    .A2(_11459_),
    .ZN(_12658_));
 AND2_X1 _22349_ (.A1(_11533_),
    .A2(_11371_),
    .ZN(_12659_));
 NOR4_X1 _22350_ (.A1(_12656_),
    .A2(_12657_),
    .A3(_12658_),
    .A4(_12659_),
    .ZN(_12660_));
 INV_X1 _22351_ (.A(_11529_),
    .ZN(_12661_));
 NAND2_X1 _22352_ (.A1(_11431_),
    .A2(_11461_),
    .ZN(_12662_));
 AND4_X1 _22353_ (.A1(_11494_),
    .A2(_12661_),
    .A3(_12662_),
    .A4(_11468_),
    .ZN(_12663_));
 NOR2_X1 _22354_ (.A1(_11355_),
    .A2(_11418_),
    .ZN(_12664_));
 AND2_X1 _22355_ (.A1(_11366_),
    .A2(_12664_),
    .ZN(_12665_));
 INV_X1 _22356_ (.A(_12665_),
    .ZN(_12666_));
 AND2_X1 _22357_ (.A1(_11477_),
    .A2(_12296_),
    .ZN(_12667_));
 INV_X1 _22358_ (.A(_12667_),
    .ZN(_12668_));
 AND2_X1 _22359_ (.A1(_11352_),
    .A2(_12322_),
    .ZN(_12669_));
 INV_X1 _22360_ (.A(_12669_),
    .ZN(_12670_));
 NAND2_X1 _22361_ (.A1(_11400_),
    .A2(_11318_),
    .ZN(_12671_));
 AND4_X1 _22362_ (.A1(_12666_),
    .A2(_12668_),
    .A3(_12670_),
    .A4(_12671_),
    .ZN(_12672_));
 AND4_X1 _22363_ (.A1(_12655_),
    .A2(_12660_),
    .A3(_12663_),
    .A4(_12672_),
    .ZN(_12673_));
 NAND2_X1 _22364_ (.A1(_12375_),
    .A2(_11406_),
    .ZN(_12674_));
 NAND4_X1 _22365_ (.A1(_11323_),
    .A2(_12674_),
    .A3(_12370_),
    .A4(_12307_),
    .ZN(_12675_));
 OAI22_X1 _22366_ (.A1(_11434_),
    .A2(_12374_),
    .B1(_12296_),
    .B2(_11489_),
    .ZN(_12676_));
 NAND3_X1 _22367_ (.A1(_12366_),
    .A2(_11408_),
    .A3(_11356_),
    .ZN(_12677_));
 NAND2_X1 _22368_ (.A1(_12338_),
    .A2(_11406_),
    .ZN(_12678_));
 NAND4_X1 _22369_ (.A1(_12676_),
    .A2(_12294_),
    .A3(_12677_),
    .A4(_12678_),
    .ZN(_12679_));
 NOR4_X1 _22370_ (.A1(_12675_),
    .A2(_12679_),
    .A3(_11348_),
    .A4(_11471_),
    .ZN(_12680_));
 AND2_X1 _22371_ (.A1(_11330_),
    .A2(_11429_),
    .ZN(_12681_));
 NOR2_X1 _22372_ (.A1(_11476_),
    .A2(_12681_),
    .ZN(_12682_));
 OAI21_X1 _22373_ (.A(_11497_),
    .B1(_11400_),
    .B2(_11420_),
    .ZN(_12683_));
 OAI21_X1 _22374_ (.A(_11497_),
    .B1(_12296_),
    .B2(_11525_),
    .ZN(_12684_));
 AND2_X1 _22375_ (.A1(_12683_),
    .A2(_12684_),
    .ZN(_12685_));
 AND4_X1 _22376_ (.A1(_11388_),
    .A2(_11334_),
    .A3(_11351_),
    .A4(_11365_),
    .ZN(_12686_));
 NOR2_X1 _22377_ (.A1(_11430_),
    .A2(_12686_),
    .ZN(_12687_));
 OAI21_X1 _22378_ (.A(_11460_),
    .B1(_11444_),
    .B2(_11456_),
    .ZN(_12688_));
 AND4_X1 _22379_ (.A1(_12682_),
    .A2(_12685_),
    .A3(_12687_),
    .A4(_12688_),
    .ZN(_12689_));
 NOR2_X1 _22380_ (.A1(_11469_),
    .A2(_11418_),
    .ZN(_12690_));
 AND2_X1 _22381_ (.A1(_11352_),
    .A2(_12690_),
    .ZN(_12691_));
 INV_X1 _22382_ (.A(_12691_),
    .ZN(_12692_));
 AOI22_X1 _22383_ (.A1(_11518_),
    .A2(_12366_),
    .B1(_11481_),
    .B2(_11437_),
    .ZN(_12693_));
 INV_X1 _22384_ (.A(_11353_),
    .ZN(_12694_));
 OAI211_X1 _22385_ (.A(_12692_),
    .B(_12693_),
    .C1(_12318_),
    .C2(_12694_),
    .ZN(_12695_));
 AOI22_X1 _22386_ (.A1(_11403_),
    .A2(_11456_),
    .B1(_11398_),
    .B2(_11431_),
    .ZN(_12696_));
 INV_X1 _22387_ (.A(_11405_),
    .ZN(_12697_));
 OAI221_X1 _22388_ (.A(_12696_),
    .B1(_11441_),
    .B2(_12697_),
    .C1(_11539_),
    .C2(_12345_),
    .ZN(_12698_));
 AOI22_X1 _22389_ (.A1(_11344_),
    .A2(_12374_),
    .B1(_12338_),
    .B2(_11536_),
    .ZN(_12699_));
 NAND2_X1 _22390_ (.A1(_11481_),
    .A2(_12690_),
    .ZN(_12700_));
 NAND2_X1 _22391_ (.A1(_11427_),
    .A2(_11490_),
    .ZN(_12701_));
 NAND3_X1 _22392_ (.A1(_12699_),
    .A2(_12700_),
    .A3(_12701_),
    .ZN(_12702_));
 AOI22_X1 _22393_ (.A1(_11493_),
    .A2(_11414_),
    .B1(_11511_),
    .B2(_11536_),
    .ZN(_12703_));
 NAND2_X1 _22394_ (.A1(_11353_),
    .A2(_12338_),
    .ZN(_12704_));
 NAND3_X1 _22395_ (.A1(_11415_),
    .A2(_11338_),
    .A3(_11359_),
    .ZN(_12705_));
 NAND3_X1 _22396_ (.A1(_12703_),
    .A2(_12704_),
    .A3(_12705_),
    .ZN(_12706_));
 NOR4_X1 _22397_ (.A1(_12695_),
    .A2(_12698_),
    .A3(_12702_),
    .A4(_12706_),
    .ZN(_12707_));
 NAND4_X1 _22398_ (.A1(_12673_),
    .A2(_12680_),
    .A3(_12689_),
    .A4(_12707_),
    .ZN(_12708_));
 OAI21_X1 _22399_ (.A(_11483_),
    .B1(_11344_),
    .B2(_11456_),
    .ZN(_12709_));
 NAND4_X1 _22400_ (.A1(_11381_),
    .A2(_11389_),
    .A3(_11385_),
    .A4(_11435_),
    .ZN(_12710_));
 NAND4_X1 _22401_ (.A1(_11483_),
    .A2(_11396_),
    .A3(_11408_),
    .A4(_11388_),
    .ZN(_12711_));
 NAND3_X1 _22402_ (.A1(_12709_),
    .A2(_12710_),
    .A3(_12711_),
    .ZN(_12712_));
 AND2_X1 _22403_ (.A1(_11481_),
    .A2(_11518_),
    .ZN(_12713_));
 INV_X1 _22404_ (.A(_12713_),
    .ZN(_12714_));
 INV_X1 _22405_ (.A(_11518_),
    .ZN(_12715_));
 OAI221_X1 _22406_ (.A(_12714_),
    .B1(_12313_),
    .B2(_11524_),
    .C1(_12715_),
    .C2(_11440_),
    .ZN(_12716_));
 AND2_X1 _22407_ (.A1(_11507_),
    .A2(_11407_),
    .ZN(_12717_));
 AOI22_X1 _22408_ (.A1(_12717_),
    .A2(_11415_),
    .B1(_11542_),
    .B2(_12374_),
    .ZN(_12718_));
 NAND2_X1 _22409_ (.A1(_12664_),
    .A2(_11487_),
    .ZN(_12719_));
 AND2_X1 _22410_ (.A1(_12719_),
    .A2(_12316_),
    .ZN(_12720_));
 OAI21_X1 _22411_ (.A(_11522_),
    .B1(_11410_),
    .B2(_11371_),
    .ZN(_12721_));
 NAND3_X1 _22412_ (.A1(_12718_),
    .A2(_12720_),
    .A3(_12721_),
    .ZN(_12722_));
 OAI21_X1 _22413_ (.A(_11481_),
    .B1(_12338_),
    .B2(_12296_),
    .ZN(_12723_));
 INV_X1 _22414_ (.A(_11370_),
    .ZN(_12724_));
 OAI221_X1 _22415_ (.A(_12723_),
    .B1(_12329_),
    .B2(_12724_),
    .C1(_11378_),
    .C2(_12694_),
    .ZN(_12725_));
 OR4_X1 _22416_ (.A1(_12712_),
    .A2(_12716_),
    .A3(_12722_),
    .A4(_12725_),
    .ZN(_12726_));
 NOR2_X2 _22417_ (.A1(_12708_),
    .A2(_12726_),
    .ZN(_12727_));
 XNOR2_X1 _22418_ (.A(_12651_),
    .B(_12727_),
    .ZN(_12728_));
 AND2_X1 _22419_ (.A1(_12019_),
    .A2(_12003_),
    .ZN(_12729_));
 INV_X1 _22420_ (.A(_12729_),
    .ZN(_12730_));
 NAND2_X1 _22421_ (.A1(_11964_),
    .A2(_11926_),
    .ZN(_12731_));
 AOI22_X1 _22422_ (.A1(_11959_),
    .A2(_12048_),
    .B1(_12092_),
    .B2(_11985_),
    .ZN(_12732_));
 AND4_X1 _22423_ (.A1(_12420_),
    .A2(_12730_),
    .A3(_12731_),
    .A4(_12732_),
    .ZN(_12733_));
 AOI22_X1 _22424_ (.A1(_12090_),
    .A2(_12391_),
    .B1(_12024_),
    .B2(_12089_),
    .ZN(_12734_));
 AOI221_X4 _22425_ (.A(_11949_),
    .B1(_11925_),
    .B2(_11937_),
    .C1(_12449_),
    .C2(_12088_),
    .ZN(_12735_));
 AND4_X1 _22426_ (.A1(_12404_),
    .A2(_12733_),
    .A3(_12734_),
    .A4(_12735_),
    .ZN(_12736_));
 BUF_X2 _22427_ (.A(_11962_),
    .Z(_12737_));
 NAND2_X1 _22428_ (.A1(_12000_),
    .A2(_12737_),
    .ZN(_12738_));
 NAND2_X1 _22429_ (.A1(_12006_),
    .A2(_12080_),
    .ZN(_12739_));
 INV_X1 _22430_ (.A(_12006_),
    .ZN(_12740_));
 OAI211_X1 _22431_ (.A(_12738_),
    .B(_12739_),
    .C1(_12740_),
    .C2(_11991_),
    .ZN(_12741_));
 INV_X1 _22432_ (.A(_12088_),
    .ZN(_12742_));
 INV_X1 _22433_ (.A(_12003_),
    .ZN(_12743_));
 AOI21_X1 _22434_ (.A(_12742_),
    .B1(_12426_),
    .B2(_12743_),
    .ZN(_12744_));
 AND2_X1 _22435_ (.A1(_12068_),
    .A2(_12048_),
    .ZN(_12745_));
 OR3_X1 _22436_ (.A1(_12741_),
    .A2(_12744_),
    .A3(_12745_),
    .ZN(_12746_));
 NOR2_X1 _22437_ (.A1(_11980_),
    .A2(_11907_),
    .ZN(_12747_));
 OAI21_X1 _22438_ (.A(_11914_),
    .B1(_12481_),
    .B2(_12747_),
    .ZN(_12748_));
 NAND3_X1 _22439_ (.A1(_12455_),
    .A2(_11911_),
    .A3(_12018_),
    .ZN(_12749_));
 NAND4_X1 _22440_ (.A1(_12021_),
    .A2(_12060_),
    .A3(_12043_),
    .A4(_12749_),
    .ZN(_12750_));
 NAND3_X1 _22441_ (.A1(_12064_),
    .A2(_11932_),
    .A3(_11948_),
    .ZN(_12751_));
 NAND2_X1 _22442_ (.A1(_12410_),
    .A2(_11943_),
    .ZN(_12752_));
 INV_X2 _22443_ (.A(_11942_),
    .ZN(_12753_));
 OAI211_X1 _22444_ (.A(_12751_),
    .B(_12752_),
    .C1(_12387_),
    .C2(_12753_),
    .ZN(_12754_));
 NOR4_X1 _22445_ (.A1(_12746_),
    .A2(_12748_),
    .A3(_12750_),
    .A4(_12754_),
    .ZN(_12755_));
 INV_X1 _22446_ (.A(_12092_),
    .ZN(_12756_));
 NOR2_X1 _22447_ (.A1(_12756_),
    .A2(_12398_),
    .ZN(_12757_));
 NOR2_X1 _22448_ (.A1(_12742_),
    .A2(_12416_),
    .ZN(_12758_));
 AND3_X1 _22449_ (.A1(_12030_),
    .A2(_12397_),
    .A3(_11944_),
    .ZN(_12759_));
 AND2_X1 _22450_ (.A1(_12030_),
    .A2(_12011_),
    .ZN(_12760_));
 NOR4_X1 _22451_ (.A1(_12757_),
    .A2(_12758_),
    .A3(_12759_),
    .A4(_12760_),
    .ZN(_12761_));
 BUF_X2 _22452_ (.A(_11887_),
    .Z(_12762_));
 BUF_X2 _22453_ (.A(_12048_),
    .Z(_12763_));
 AOI22_X1 _22454_ (.A1(_12762_),
    .A2(_12763_),
    .B1(_12737_),
    .B2(_12489_),
    .ZN(_12764_));
 NAND3_X1 _22455_ (.A1(_11894_),
    .A2(_11977_),
    .A3(_11979_),
    .ZN(_12765_));
 NAND2_X1 _22456_ (.A1(_12737_),
    .A2(_12762_),
    .ZN(_12766_));
 AND4_X1 _22457_ (.A1(_12056_),
    .A2(_12764_),
    .A3(_12765_),
    .A4(_12766_),
    .ZN(_12767_));
 AND4_X1 _22458_ (.A1(_12736_),
    .A2(_12755_),
    .A3(_12761_),
    .A4(_12767_),
    .ZN(_12768_));
 NAND3_X1 _22459_ (.A1(_11898_),
    .A2(_11977_),
    .A3(_11912_),
    .ZN(_12769_));
 AND4_X1 _22460_ (.A1(_11893_),
    .A2(_11978_),
    .A3(_11920_),
    .A4(_11941_),
    .ZN(_12770_));
 NOR2_X1 _22461_ (.A1(_12453_),
    .A2(_12770_),
    .ZN(_12771_));
 NAND4_X1 _22462_ (.A1(_11977_),
    .A2(_11945_),
    .A3(_11912_),
    .A4(_11955_),
    .ZN(_12772_));
 NAND3_X1 _22463_ (.A1(_11882_),
    .A2(_11977_),
    .A3(_11912_),
    .ZN(_12773_));
 AND4_X1 _22464_ (.A1(_12769_),
    .A2(_12771_),
    .A3(_12772_),
    .A4(_12773_),
    .ZN(_12774_));
 AND2_X1 _22465_ (.A1(_12009_),
    .A2(_12401_),
    .ZN(_12775_));
 AND2_X1 _22466_ (.A1(_11974_),
    .A2(_11994_),
    .ZN(_12776_));
 AOI211_X1 _22467_ (.A(_12775_),
    .B(_12776_),
    .C1(_12489_),
    .C2(_12412_),
    .ZN(_12777_));
 INV_X1 _22468_ (.A(_12498_),
    .ZN(_12778_));
 NAND2_X1 _22469_ (.A1(_11974_),
    .A2(_11937_),
    .ZN(_12779_));
 AND2_X1 _22470_ (.A1(_11944_),
    .A2(_11932_),
    .ZN(_12780_));
 INV_X1 _22471_ (.A(_12780_),
    .ZN(_12781_));
 OAI21_X1 _22472_ (.A(_12779_),
    .B1(_12044_),
    .B2(_12781_),
    .ZN(_12782_));
 AND2_X1 _22473_ (.A1(_12068_),
    .A2(_11994_),
    .ZN(_12783_));
 AND3_X1 _22474_ (.A1(_12762_),
    .A2(_11933_),
    .A3(_12010_),
    .ZN(_12784_));
 AND3_X1 _22475_ (.A1(_12455_),
    .A2(_11924_),
    .A3(_11979_),
    .ZN(_12785_));
 NOR4_X1 _22476_ (.A1(_12782_),
    .A2(_12783_),
    .A3(_12784_),
    .A4(_12785_),
    .ZN(_12786_));
 NAND4_X1 _22477_ (.A1(_12774_),
    .A2(_12777_),
    .A3(_12778_),
    .A4(_12786_),
    .ZN(_12787_));
 AND2_X1 _22478_ (.A1(_12078_),
    .A2(_12010_),
    .ZN(_12788_));
 AOI21_X1 _22479_ (.A(_12079_),
    .B1(_12395_),
    .B2(_12075_),
    .ZN(_12789_));
 NOR2_X1 _22480_ (.A1(_12033_),
    .A2(_11987_),
    .ZN(_12790_));
 AOI21_X1 _22481_ (.A(_12069_),
    .B1(_12790_),
    .B2(_12747_),
    .ZN(_12791_));
 NOR2_X1 _22482_ (.A1(_12079_),
    .A2(_12398_),
    .ZN(_12792_));
 OR4_X1 _22483_ (.A1(_12788_),
    .A2(_12789_),
    .A3(_12791_),
    .A4(_12792_),
    .ZN(_12793_));
 AND2_X1 _22484_ (.A1(_12417_),
    .A2(_12063_),
    .ZN(_12794_));
 INV_X1 _22485_ (.A(_12794_),
    .ZN(_12795_));
 OAI21_X1 _22486_ (.A(_11993_),
    .B1(_11970_),
    .B2(_11980_),
    .ZN(_12796_));
 OAI21_X1 _22487_ (.A(_12440_),
    .B1(_11970_),
    .B2(_12034_),
    .ZN(_12797_));
 OAI21_X1 _22488_ (.A(_12423_),
    .B1(_12090_),
    .B2(_12780_),
    .ZN(_12798_));
 NAND4_X1 _22489_ (.A1(_12795_),
    .A2(_12796_),
    .A3(_12797_),
    .A4(_12798_),
    .ZN(_12799_));
 OAI21_X1 _22490_ (.A(_11943_),
    .B1(_11989_),
    .B2(_12449_),
    .ZN(_12800_));
 AND2_X1 _22491_ (.A1(_11973_),
    .A2(_11904_),
    .ZN(_12801_));
 INV_X1 _22492_ (.A(_12801_),
    .ZN(_12802_));
 NAND2_X1 _22493_ (.A1(_12009_),
    .A2(_12438_),
    .ZN(_12803_));
 OAI21_X1 _22494_ (.A(_12461_),
    .B1(_12394_),
    .B2(_12425_),
    .ZN(_12804_));
 NAND4_X1 _22495_ (.A1(_12800_),
    .A2(_12802_),
    .A3(_12803_),
    .A4(_12804_),
    .ZN(_12805_));
 NOR4_X1 _22496_ (.A1(_12787_),
    .A2(_12793_),
    .A3(_12799_),
    .A4(_12805_),
    .ZN(_12806_));
 NAND2_X2 _22497_ (.A1(_12768_),
    .A2(_12806_),
    .ZN(_12807_));
 XNOR2_X1 _22498_ (.A(_12181_),
    .B(_12807_),
    .ZN(_12808_));
 XNOR2_X1 _22499_ (.A(_12728_),
    .B(_12808_),
    .ZN(_12809_));
 XNOR2_X1 _22500_ (.A(_12809_),
    .B(_17185_),
    .ZN(_12810_));
 MUX2_X1 _22501_ (.A(_12503_),
    .B(_12810_),
    .S(_11084_),
    .Z(_00718_));
 XOR2_X1 _22502_ (.A(_17188_),
    .B(_16991_),
    .Z(_12811_));
 NAND4_X1 _22503_ (.A1(_11193_),
    .A2(_11143_),
    .A3(_11239_),
    .A4(_11142_),
    .ZN(_12812_));
 INV_X1 _22504_ (.A(_11206_),
    .ZN(_12813_));
 NAND2_X1 _22505_ (.A1(_11205_),
    .A2(_11281_),
    .ZN(_12814_));
 OAI21_X1 _22506_ (.A(_11205_),
    .B1(_11248_),
    .B2(_11180_),
    .ZN(_12815_));
 NAND3_X1 _22507_ (.A1(_11215_),
    .A2(_11170_),
    .A3(_12182_),
    .ZN(_12816_));
 AND4_X1 _22508_ (.A1(_12813_),
    .A2(_12814_),
    .A3(_12815_),
    .A4(_12816_),
    .ZN(_12817_));
 OAI211_X1 _22509_ (.A(_11175_),
    .B(_11194_),
    .C1(_11125_),
    .C2(_11155_),
    .ZN(_12818_));
 AND4_X1 _22510_ (.A1(_11115_),
    .A2(_11114_),
    .A3(_11170_),
    .A4(_11135_),
    .ZN(_12819_));
 AOI221_X4 _22511_ (.A(_12819_),
    .B1(_11171_),
    .B2(_11121_),
    .C1(_12247_),
    .C2(_11124_),
    .ZN(_12820_));
 AND4_X1 _22512_ (.A1(_12812_),
    .A2(_12817_),
    .A3(_12818_),
    .A4(_12820_),
    .ZN(_12821_));
 AND2_X1 _22513_ (.A1(_12186_),
    .A2(_16738_),
    .ZN(_12822_));
 OAI21_X1 _22514_ (.A(_11129_),
    .B1(_11128_),
    .B2(_12822_),
    .ZN(_12823_));
 NAND4_X1 _22515_ (.A1(_11129_),
    .A2(_11184_),
    .A3(_11186_),
    .A4(_11099_),
    .ZN(_12824_));
 AND2_X1 _22516_ (.A1(_12824_),
    .A2(_11106_),
    .ZN(_12825_));
 OAI21_X1 _22517_ (.A(_11092_),
    .B1(_11177_),
    .B2(_11190_),
    .ZN(_12826_));
 OAI21_X1 _22518_ (.A(_11092_),
    .B1(_12233_),
    .B2(_11162_),
    .ZN(_12827_));
 AND4_X1 _22519_ (.A1(_12823_),
    .A2(_12825_),
    .A3(_12826_),
    .A4(_12827_),
    .ZN(_12828_));
 AND2_X2 _22520_ (.A1(_11125_),
    .A2(_11114_),
    .ZN(_12829_));
 AND2_X1 _22521_ (.A1(_11126_),
    .A2(_11124_),
    .ZN(_12830_));
 OAI21_X1 _22522_ (.A(_11137_),
    .B1(_12829_),
    .B2(_12830_),
    .ZN(_12831_));
 OAI21_X1 _22523_ (.A(_11136_),
    .B1(_11248_),
    .B2(_11181_),
    .ZN(_12832_));
 NAND3_X1 _22524_ (.A1(_12831_),
    .A2(_12212_),
    .A3(_12832_),
    .ZN(_12833_));
 NAND2_X1 _22525_ (.A1(_11148_),
    .A2(_11304_),
    .ZN(_12834_));
 OAI211_X1 _22526_ (.A(_12223_),
    .B(_12834_),
    .C1(_12224_),
    .C2(_12198_),
    .ZN(_12835_));
 NAND2_X1 _22527_ (.A1(_11148_),
    .A2(_11133_),
    .ZN(_12836_));
 NAND2_X1 _22528_ (.A1(_11148_),
    .A2(_11105_),
    .ZN(_12837_));
 NAND2_X1 _22529_ (.A1(_12836_),
    .A2(_12837_),
    .ZN(_12838_));
 NOR3_X1 _22530_ (.A1(_12833_),
    .A2(_12835_),
    .A3(_12838_),
    .ZN(_12839_));
 AOI21_X1 _22531_ (.A(_11214_),
    .B1(_12623_),
    .B2(_12192_),
    .ZN(_12840_));
 AND3_X1 _22532_ (.A1(_11230_),
    .A2(_11203_),
    .A3(_11191_),
    .ZN(_12841_));
 AND2_X1 _22533_ (.A1(_11213_),
    .A2(_11127_),
    .ZN(_12842_));
 AND2_X1 _22534_ (.A1(_11215_),
    .A2(_11191_),
    .ZN(_12843_));
 NOR4_X1 _22535_ (.A1(_12840_),
    .A2(_12841_),
    .A3(_12842_),
    .A4(_12843_),
    .ZN(_12844_));
 NAND4_X1 _22536_ (.A1(_12821_),
    .A2(_12828_),
    .A3(_12839_),
    .A4(_12844_),
    .ZN(_12845_));
 AOI21_X1 _22537_ (.A(_12607_),
    .B1(_12618_),
    .B2(_12219_),
    .ZN(_12846_));
 AND4_X1 _22538_ (.A1(_11231_),
    .A2(_11098_),
    .A3(_11189_),
    .A4(_11135_),
    .ZN(_12847_));
 OR3_X1 _22539_ (.A1(_12846_),
    .A2(_12608_),
    .A3(_12847_),
    .ZN(_12848_));
 AND2_X1 _22540_ (.A1(_12580_),
    .A2(_11252_),
    .ZN(_12849_));
 OAI21_X1 _22541_ (.A(_12605_),
    .B1(_12266_),
    .B2(_12192_),
    .ZN(_12850_));
 NOR4_X1 _22542_ (.A1(_12848_),
    .A2(_12849_),
    .A3(_12264_),
    .A4(_12850_),
    .ZN(_12851_));
 OAI21_X1 _22543_ (.A(_11285_),
    .B1(_11267_),
    .B2(_12275_),
    .ZN(_12852_));
 OAI21_X1 _22544_ (.A(_11285_),
    .B1(_12205_),
    .B2(_11282_),
    .ZN(_12853_));
 OAI21_X1 _22545_ (.A(_11274_),
    .B1(_11301_),
    .B2(_11116_),
    .ZN(_12854_));
 OAI211_X1 _22546_ (.A(_11088_),
    .B(_11288_),
    .C1(_11215_),
    .C2(_11217_),
    .ZN(_12855_));
 NAND4_X1 _22547_ (.A1(_12852_),
    .A2(_12853_),
    .A3(_12854_),
    .A4(_12855_),
    .ZN(_12856_));
 NAND2_X1 _22548_ (.A1(_12829_),
    .A2(_11297_),
    .ZN(_12857_));
 OAI211_X1 _22549_ (.A(_12857_),
    .B(_11307_),
    .C1(_12219_),
    .C2(_12208_),
    .ZN(_12858_));
 AOI21_X1 _22550_ (.A(_12208_),
    .B1(_11278_),
    .B2(_11210_),
    .ZN(_12859_));
 OAI21_X1 _22551_ (.A(_11298_),
    .B1(_12227_),
    .B2(_12208_),
    .ZN(_12860_));
 NOR4_X1 _22552_ (.A1(_12856_),
    .A2(_12858_),
    .A3(_12859_),
    .A4(_12860_),
    .ZN(_12861_));
 INV_X1 _22553_ (.A(_11264_),
    .ZN(_12862_));
 INV_X1 _22554_ (.A(_11159_),
    .ZN(_12863_));
 NAND2_X1 _22555_ (.A1(_12227_),
    .A2(_12863_),
    .ZN(_12864_));
 INV_X1 _22556_ (.A(_12864_),
    .ZN(_12865_));
 AOI21_X1 _22557_ (.A(_12862_),
    .B1(_12865_),
    .B2(_12623_),
    .ZN(_12866_));
 AND2_X1 _22558_ (.A1(_11116_),
    .A2(_11264_),
    .ZN(_12867_));
 OAI21_X1 _22559_ (.A(_11291_),
    .B1(_11138_),
    .B2(_11217_),
    .ZN(_12868_));
 OAI211_X1 _22560_ (.A(_11291_),
    .B(_11141_),
    .C1(_11109_),
    .C2(_11095_),
    .ZN(_12869_));
 OAI21_X1 _22561_ (.A(_11291_),
    .B1(_11105_),
    .B2(_11110_),
    .ZN(_12870_));
 NAND4_X1 _22562_ (.A1(_11099_),
    .A2(_11189_),
    .A3(_11288_),
    .A4(_11135_),
    .ZN(_12871_));
 NAND4_X1 _22563_ (.A1(_12868_),
    .A2(_12869_),
    .A3(_12870_),
    .A4(_12871_),
    .ZN(_12872_));
 NOR4_X1 _22564_ (.A1(_12866_),
    .A2(_12579_),
    .A3(_12867_),
    .A4(_12872_),
    .ZN(_12873_));
 OAI21_X1 _22565_ (.A(_11247_),
    .B1(_11127_),
    .B2(_11235_),
    .ZN(_12874_));
 OAI21_X1 _22566_ (.A(_12874_),
    .B1(_12616_),
    .B2(_12257_),
    .ZN(_12875_));
 OAI211_X1 _22567_ (.A(_11088_),
    .B(_11237_),
    .C1(_11163_),
    .C2(_12187_),
    .ZN(_12876_));
 NAND2_X1 _22568_ (.A1(_11259_),
    .A2(_12226_),
    .ZN(_12877_));
 NAND4_X1 _22569_ (.A1(_12876_),
    .A2(_11260_),
    .A3(_12877_),
    .A4(_12279_),
    .ZN(_12878_));
 AND4_X1 _22570_ (.A1(_11095_),
    .A2(_11237_),
    .A3(_11153_),
    .A4(_11102_),
    .ZN(_12879_));
 AOI21_X1 _22571_ (.A(_12257_),
    .B1(_12589_),
    .B2(_12863_),
    .ZN(_12880_));
 NOR4_X1 _22572_ (.A1(_12875_),
    .A2(_12878_),
    .A3(_12879_),
    .A4(_12880_),
    .ZN(_12881_));
 NAND4_X1 _22573_ (.A1(_12851_),
    .A2(_12861_),
    .A3(_12873_),
    .A4(_12881_),
    .ZN(_12882_));
 NOR2_X2 _22574_ (.A1(_12845_),
    .A2(_12882_),
    .ZN(_12883_));
 AND4_X1 _22575_ (.A1(_11620_),
    .A2(_11637_),
    .A3(_11710_),
    .A4(_11588_),
    .ZN(_12884_));
 AND4_X1 _22576_ (.A1(_11642_),
    .A2(_11620_),
    .A3(_11637_),
    .A4(_11588_),
    .ZN(_12885_));
 AOI211_X1 _22577_ (.A(_12884_),
    .B(_12885_),
    .C1(_11698_),
    .C2(_11667_),
    .ZN(_12886_));
 AOI21_X1 _22578_ (.A(_12544_),
    .B1(_11780_),
    .B2(_11845_),
    .ZN(_12887_));
 AND2_X1 _22579_ (.A1(_11664_),
    .A2(_11833_),
    .ZN(_12888_));
 NOR4_X1 _22580_ (.A1(_12887_),
    .A2(_11665_),
    .A3(_12163_),
    .A4(_12888_),
    .ZN(_12889_));
 NAND4_X1 _22581_ (.A1(_11667_),
    .A2(_11571_),
    .A3(_11671_),
    .A4(_11788_),
    .ZN(_12890_));
 OAI21_X1 _22582_ (.A(_11667_),
    .B1(_12506_),
    .B2(_11644_),
    .ZN(_12891_));
 AND4_X1 _22583_ (.A1(_12886_),
    .A2(_12889_),
    .A3(_12890_),
    .A4(_12891_),
    .ZN(_12892_));
 OAI211_X1 _22584_ (.A(_11764_),
    .B(_11570_),
    .C1(_11567_),
    .C2(_11642_),
    .ZN(_12893_));
 OAI211_X1 _22585_ (.A(_11764_),
    .B(_11620_),
    .C1(_11710_),
    .C2(_11583_),
    .ZN(_12894_));
 OAI21_X1 _22586_ (.A(_11764_),
    .B1(_11757_),
    .B2(_11687_),
    .ZN(_12895_));
 AND4_X1 _22587_ (.A1(_11771_),
    .A2(_12893_),
    .A3(_12894_),
    .A4(_12895_),
    .ZN(_12896_));
 AND2_X1 _22588_ (.A1(_11755_),
    .A2(_11621_),
    .ZN(_12897_));
 AND3_X1 _22589_ (.A1(_11694_),
    .A2(_11731_),
    .A3(_11616_),
    .ZN(_12898_));
 AND3_X1 _22590_ (.A1(_11627_),
    .A2(_11731_),
    .A3(_11616_),
    .ZN(_12899_));
 NOR4_X1 _22591_ (.A1(_12897_),
    .A2(_12898_),
    .A3(_12118_),
    .A4(_12899_),
    .ZN(_12900_));
 OAI21_X1 _22592_ (.A(_11756_),
    .B1(_11737_),
    .B2(_11587_),
    .ZN(_12901_));
 OAI211_X1 _22593_ (.A(_11732_),
    .B(_11659_),
    .C1(_11674_),
    .C2(_11643_),
    .ZN(_12902_));
 AND4_X1 _22594_ (.A1(_12896_),
    .A2(_12900_),
    .A3(_12901_),
    .A4(_12902_),
    .ZN(_12903_));
 NAND3_X1 _22595_ (.A1(_11649_),
    .A2(_11734_),
    .A3(_11788_),
    .ZN(_12904_));
 NAND4_X1 _22596_ (.A1(_11795_),
    .A2(_12570_),
    .A3(_12567_),
    .A4(_12904_),
    .ZN(_12905_));
 AOI21_X1 _22597_ (.A(_11747_),
    .B1(_11811_),
    .B2(_11691_),
    .ZN(_12906_));
 NAND4_X1 _22598_ (.A1(_11731_),
    .A2(_11583_),
    .A3(_11592_),
    .A4(_11552_),
    .ZN(_12907_));
 NAND4_X1 _22599_ (.A1(_11672_),
    .A2(_11731_),
    .A3(_11710_),
    .A4(_11552_),
    .ZN(_12908_));
 OAI211_X1 _22600_ (.A(_12907_),
    .B(_12908_),
    .C1(_11747_),
    .C2(_11595_),
    .ZN(_12909_));
 AOI21_X1 _22601_ (.A(_11747_),
    .B1(_11746_),
    .B2(_11840_),
    .ZN(_12910_));
 NOR4_X1 _22602_ (.A1(_12905_),
    .A2(_12906_),
    .A3(_12909_),
    .A4(_12910_),
    .ZN(_12911_));
 OAI21_X1 _22603_ (.A(_11656_),
    .B1(_12171_),
    .B2(_11768_),
    .ZN(_12912_));
 NAND4_X1 _22604_ (.A1(_11672_),
    .A2(_11646_),
    .A3(_11710_),
    .A4(_11572_),
    .ZN(_12913_));
 NAND3_X1 _22605_ (.A1(_12912_),
    .A2(_12554_),
    .A3(_12913_),
    .ZN(_12914_));
 AND2_X1 _22606_ (.A1(_11639_),
    .A2(_11705_),
    .ZN(_12915_));
 INV_X1 _22607_ (.A(_11598_),
    .ZN(_12916_));
 AOI21_X1 _22608_ (.A(_11783_),
    .B1(_11718_),
    .B2(_12916_),
    .ZN(_12917_));
 NOR4_X1 _22609_ (.A1(_12914_),
    .A2(_11782_),
    .A3(_12915_),
    .A4(_12917_),
    .ZN(_12918_));
 NAND4_X1 _22610_ (.A1(_12892_),
    .A2(_12903_),
    .A3(_12911_),
    .A4(_12918_),
    .ZN(_12919_));
 NAND2_X1 _22611_ (.A1(_11607_),
    .A2(_11705_),
    .ZN(_12920_));
 AOI21_X1 _22612_ (.A(_11847_),
    .B1(_11718_),
    .B2(_11758_),
    .ZN(_12921_));
 AOI21_X1 _22613_ (.A(_11847_),
    .B1(_11778_),
    .B2(_11873_),
    .ZN(_12922_));
 NOR3_X1 _22614_ (.A1(_12921_),
    .A2(_12922_),
    .A3(_12145_),
    .ZN(_12923_));
 OAI21_X1 _22615_ (.A(_11607_),
    .B1(_11737_),
    .B2(_11768_),
    .ZN(_12924_));
 OAI21_X1 _22616_ (.A(_11603_),
    .B1(_11598_),
    .B2(_11612_),
    .ZN(_12925_));
 AND4_X1 _22617_ (.A1(_12920_),
    .A2(_12923_),
    .A3(_12924_),
    .A4(_12925_),
    .ZN(_12926_));
 AND3_X1 _22618_ (.A1(_11713_),
    .A2(_11626_),
    .A3(_11620_),
    .ZN(_12927_));
 AOI211_X1 _22619_ (.A(_12927_),
    .B(_12131_),
    .C1(_11713_),
    .C2(_11698_),
    .ZN(_12928_));
 AND2_X1 _22620_ (.A1(_11679_),
    .A2(_11674_),
    .ZN(_12929_));
 AND2_X1 _22621_ (.A1(_11689_),
    .A2(_11679_),
    .ZN(_12930_));
 AOI211_X1 _22622_ (.A(_12929_),
    .B(_12930_),
    .C1(_11587_),
    .C2(_11680_),
    .ZN(_12931_));
 AOI21_X1 _22623_ (.A(_11717_),
    .B1(_11860_),
    .B2(_12108_),
    .ZN(_12932_));
 AOI21_X1 _22624_ (.A(_12932_),
    .B1(_11587_),
    .B2(_11713_),
    .ZN(_12933_));
 AND2_X1 _22625_ (.A1(_11679_),
    .A2(_11621_),
    .ZN(_12934_));
 AND2_X1 _22626_ (.A1(_11679_),
    .A2(_11669_),
    .ZN(_12935_));
 NOR2_X1 _22627_ (.A1(_12934_),
    .A2(_12935_),
    .ZN(_12936_));
 AND4_X1 _22628_ (.A1(_12928_),
    .A2(_12931_),
    .A3(_12933_),
    .A4(_12936_),
    .ZN(_12937_));
 AND2_X1 _22629_ (.A1(_11570_),
    .A2(_11824_),
    .ZN(_12938_));
 OAI21_X1 _22630_ (.A(_11581_),
    .B1(_12506_),
    .B2(_12938_),
    .ZN(_12939_));
 OAI21_X1 _22631_ (.A(_11581_),
    .B1(_11685_),
    .B2(_11612_),
    .ZN(_12940_));
 OAI211_X1 _22632_ (.A(_11566_),
    .B(_11616_),
    .C1(_12506_),
    .C2(_11643_),
    .ZN(_12941_));
 NAND2_X1 _22633_ (.A1(_11617_),
    .A2(_11608_),
    .ZN(_12942_));
 AND2_X1 _22634_ (.A1(_12941_),
    .A2(_12942_),
    .ZN(_12943_));
 OAI21_X1 _22635_ (.A(_12149_),
    .B1(_11749_),
    .B2(_12150_),
    .ZN(_12944_));
 AND4_X1 _22636_ (.A1(_12939_),
    .A2(_12940_),
    .A3(_12943_),
    .A4(_12944_),
    .ZN(_12945_));
 NAND3_X1 _22637_ (.A1(_11627_),
    .A2(_11695_),
    .A3(_11616_),
    .ZN(_12946_));
 OAI21_X1 _22638_ (.A(_12946_),
    .B1(_12531_),
    .B2(_12916_),
    .ZN(_12947_));
 AND3_X1 _22639_ (.A1(_11649_),
    .A2(_11788_),
    .A3(_11696_),
    .ZN(_12948_));
 AND2_X1 _22640_ (.A1(_11674_),
    .A2(_11696_),
    .ZN(_12949_));
 NOR4_X1 _22641_ (.A1(_12947_),
    .A2(_12948_),
    .A3(_11868_),
    .A4(_12949_),
    .ZN(_12950_));
 NAND4_X1 _22642_ (.A1(_12926_),
    .A2(_12937_),
    .A3(_12945_),
    .A4(_12950_),
    .ZN(_12951_));
 NOR2_X2 _22643_ (.A1(_12919_),
    .A2(_12951_),
    .ZN(_12952_));
 XOR2_X1 _22644_ (.A(_12883_),
    .B(_12952_),
    .Z(_12953_));
 NOR2_X1 _22645_ (.A1(_11908_),
    .A2(_12477_),
    .ZN(_12954_));
 OAI21_X1 _22646_ (.A(_12954_),
    .B1(_12475_),
    .B2(_12070_),
    .ZN(_12955_));
 AOI21_X1 _22647_ (.A(_11935_),
    .B1(_11990_),
    .B2(_11938_),
    .ZN(_12956_));
 AOI21_X1 _22648_ (.A(_11935_),
    .B1(_12083_),
    .B2(_12085_),
    .ZN(_12957_));
 NOR4_X1 _22649_ (.A1(_12955_),
    .A2(_12956_),
    .A3(_11888_),
    .A4(_12957_),
    .ZN(_12958_));
 AND2_X1 _22650_ (.A1(_11974_),
    .A2(_12024_),
    .ZN(_12959_));
 AND2_X1 _22651_ (.A1(_11973_),
    .A2(_12401_),
    .ZN(_12960_));
 AND3_X1 _22652_ (.A1(_11964_),
    .A2(_11957_),
    .A3(_11978_),
    .ZN(_12961_));
 OR4_X1 _22653_ (.A1(_12959_),
    .A2(_12776_),
    .A3(_12960_),
    .A4(_12961_),
    .ZN(_12962_));
 NOR2_X1 _22654_ (.A1(_11984_),
    .A2(_12430_),
    .ZN(_12963_));
 AND2_X1 _22655_ (.A1(_11993_),
    .A2(_12414_),
    .ZN(_12964_));
 AOI211_X1 _22656_ (.A(_11916_),
    .B(_11984_),
    .C1(_11946_),
    .C2(_16785_),
    .ZN(_12965_));
 NOR4_X1 _22657_ (.A1(_12962_),
    .A2(_12963_),
    .A3(_12964_),
    .A4(_12965_),
    .ZN(_12966_));
 OAI21_X1 _22658_ (.A(_12480_),
    .B1(_12763_),
    .B2(_11929_),
    .ZN(_12967_));
 OAI21_X1 _22659_ (.A(_12480_),
    .B1(_12080_),
    .B2(_12401_),
    .ZN(_12968_));
 OAI211_X1 _22660_ (.A(_11977_),
    .B(_11912_),
    .C1(_12410_),
    .C2(_12412_),
    .ZN(_12969_));
 NAND4_X1 _22661_ (.A1(_12967_),
    .A2(_12968_),
    .A3(_12969_),
    .A4(_12773_),
    .ZN(_12970_));
 OAI21_X1 _22662_ (.A(_11943_),
    .B1(_12425_),
    .B2(_11953_),
    .ZN(_12971_));
 NAND2_X1 _22663_ (.A1(_12763_),
    .A2(_11943_),
    .ZN(_12972_));
 NAND2_X1 _22664_ (.A1(_12971_),
    .A2(_12972_),
    .ZN(_12973_));
 AOI21_X1 _22665_ (.A(_12753_),
    .B1(_12402_),
    .B2(_12013_),
    .ZN(_12974_));
 NOR3_X1 _22666_ (.A1(_12970_),
    .A2(_12973_),
    .A3(_12974_),
    .ZN(_12975_));
 INV_X1 _22667_ (.A(_12460_),
    .ZN(_12976_));
 OAI21_X1 _22668_ (.A(_12000_),
    .B1(_12003_),
    .B2(_12410_),
    .ZN(_12977_));
 OAI21_X1 _22669_ (.A(_12000_),
    .B1(_12737_),
    .B2(_11937_),
    .ZN(_12978_));
 OAI21_X1 _22670_ (.A(_12000_),
    .B1(_12763_),
    .B2(_11994_),
    .ZN(_12979_));
 AND4_X1 _22671_ (.A1(_12976_),
    .A2(_12977_),
    .A3(_12978_),
    .A4(_12979_),
    .ZN(_12980_));
 OAI211_X1 _22672_ (.A(_12009_),
    .B(_12414_),
    .C1(_11945_),
    .C2(_11946_),
    .ZN(_12981_));
 OAI21_X1 _22673_ (.A(_12009_),
    .B1(_12394_),
    .B2(_12763_),
    .ZN(_12982_));
 AND3_X1 _22674_ (.A1(_12980_),
    .A2(_12981_),
    .A3(_12982_),
    .ZN(_12983_));
 AND4_X1 _22675_ (.A1(_12958_),
    .A2(_12966_),
    .A3(_12975_),
    .A4(_12983_),
    .ZN(_12984_));
 OAI211_X1 _22676_ (.A(_12423_),
    .B(_12010_),
    .C1(_11919_),
    .C2(_11906_),
    .ZN(_12985_));
 OAI211_X1 _22677_ (.A(_12423_),
    .B(_12011_),
    .C1(_11927_),
    .C2(_11920_),
    .ZN(_12986_));
 OAI211_X1 _22678_ (.A(_12423_),
    .B(_12414_),
    .C1(_11927_),
    .C2(_11919_),
    .ZN(_12987_));
 NAND2_X1 _22679_ (.A1(_12423_),
    .A2(_12080_),
    .ZN(_12988_));
 NAND4_X1 _22680_ (.A1(_12985_),
    .A2(_12986_),
    .A3(_12987_),
    .A4(_12988_),
    .ZN(_12989_));
 NAND2_X1 _22681_ (.A1(_11953_),
    .A2(_12440_),
    .ZN(_12990_));
 NAND2_X1 _22682_ (.A1(_12053_),
    .A2(_12990_),
    .ZN(_12991_));
 NOR4_X1 _22683_ (.A1(_12989_),
    .A2(_12448_),
    .A3(_12450_),
    .A4(_12991_),
    .ZN(_12992_));
 OAI21_X1 _22684_ (.A(_12089_),
    .B1(_12399_),
    .B2(_11900_),
    .ZN(_12993_));
 OAI211_X1 _22685_ (.A(_12993_),
    .B(_12420_),
    .C1(_12085_),
    .C2(_12742_),
    .ZN(_12994_));
 NOR2_X1 _22686_ (.A1(_12756_),
    .A2(_12430_),
    .ZN(_12995_));
 AOI21_X1 _22687_ (.A(_12756_),
    .B1(_12406_),
    .B2(_11938_),
    .ZN(_12996_));
 NAND4_X1 _22688_ (.A1(_11911_),
    .A2(_12010_),
    .A3(_11920_),
    .A4(_12018_),
    .ZN(_12997_));
 NAND4_X1 _22689_ (.A1(_11911_),
    .A2(_11919_),
    .A3(_12011_),
    .A4(_12018_),
    .ZN(_12998_));
 INV_X1 _22690_ (.A(_11994_),
    .ZN(_12999_));
 OAI211_X1 _22691_ (.A(_12997_),
    .B(_12998_),
    .C1(_12756_),
    .C2(_12999_),
    .ZN(_13000_));
 NOR4_X1 _22692_ (.A1(_12994_),
    .A2(_12995_),
    .A3(_12996_),
    .A4(_13000_),
    .ZN(_13001_));
 OAI21_X1 _22693_ (.A(_12078_),
    .B1(_11898_),
    .B2(_11894_),
    .ZN(_13002_));
 OAI21_X1 _22694_ (.A(_12068_),
    .B1(_11898_),
    .B2(_12447_),
    .ZN(_13003_));
 OAI21_X1 _22695_ (.A(_12068_),
    .B1(_12763_),
    .B2(_12084_),
    .ZN(_13004_));
 OAI21_X1 _22696_ (.A(_12078_),
    .B1(_12763_),
    .B2(_12412_),
    .ZN(_13005_));
 AND4_X1 _22697_ (.A1(_13002_),
    .A2(_13003_),
    .A3(_13004_),
    .A4(_13005_),
    .ZN(_13006_));
 OAI21_X1 _22698_ (.A(_12022_),
    .B1(_12737_),
    .B2(_12447_),
    .ZN(_13007_));
 NAND2_X1 _22699_ (.A1(_12022_),
    .A2(_11964_),
    .ZN(_13008_));
 NAND4_X1 _22700_ (.A1(_12028_),
    .A2(_13007_),
    .A3(_12025_),
    .A4(_13008_),
    .ZN(_13009_));
 NAND2_X1 _22701_ (.A1(_12760_),
    .A2(_12429_),
    .ZN(_13010_));
 NAND3_X1 _22702_ (.A1(_12391_),
    .A2(_12010_),
    .A3(_11920_),
    .ZN(_13011_));
 NAND2_X1 _22703_ (.A1(_13010_),
    .A2(_13011_),
    .ZN(_13012_));
 NOR3_X1 _22704_ (.A1(_12037_),
    .A2(_11919_),
    .A3(_12416_),
    .ZN(_13013_));
 AND2_X1 _22705_ (.A1(_11882_),
    .A2(_12391_),
    .ZN(_13014_));
 NOR4_X1 _22706_ (.A1(_13009_),
    .A2(_13012_),
    .A3(_13013_),
    .A4(_13014_),
    .ZN(_13015_));
 AND4_X1 _22707_ (.A1(_12992_),
    .A2(_13001_),
    .A3(_13006_),
    .A4(_13015_),
    .ZN(_13016_));
 NAND2_X2 _22708_ (.A1(_12984_),
    .A2(_13016_),
    .ZN(_13017_));
 XNOR2_X1 _22709_ (.A(_13017_),
    .B(_12101_),
    .ZN(_13018_));
 XNOR2_X1 _22710_ (.A(_12953_),
    .B(_13018_),
    .ZN(_13019_));
 XOR2_X2 _22711_ (.A(_11877_),
    .B(_12575_),
    .Z(_13020_));
 OAI211_X1 _22712_ (.A(_11459_),
    .B(_11396_),
    .C1(_11319_),
    .C2(_11343_),
    .ZN(_13021_));
 OAI211_X1 _22713_ (.A(_11458_),
    .B(_11334_),
    .C1(_11338_),
    .C2(_11335_),
    .ZN(_13022_));
 OAI21_X1 _22714_ (.A(_11459_),
    .B1(_11442_),
    .B2(_11461_),
    .ZN(_13023_));
 AND4_X1 _22715_ (.A1(_11503_),
    .A2(_13021_),
    .A3(_13022_),
    .A4(_13023_),
    .ZN(_13024_));
 AND3_X1 _22716_ (.A1(_11424_),
    .A2(_11364_),
    .A3(_11365_),
    .ZN(_13025_));
 AOI21_X1 _22717_ (.A(_11440_),
    .B1(_11341_),
    .B2(_12298_),
    .ZN(_13026_));
 AOI211_X1 _22718_ (.A(_13025_),
    .B(_13026_),
    .C1(_11525_),
    .C2(_11366_),
    .ZN(_13027_));
 OAI21_X1 _22719_ (.A(_11434_),
    .B1(_11420_),
    .B2(_11493_),
    .ZN(_13028_));
 OAI21_X1 _22720_ (.A(_11434_),
    .B1(_11511_),
    .B2(_11437_),
    .ZN(_13029_));
 AND4_X1 _22721_ (.A1(_13024_),
    .A2(_13027_),
    .A3(_13028_),
    .A4(_13029_),
    .ZN(_13030_));
 AND2_X1 _22722_ (.A1(_11426_),
    .A2(_11327_),
    .ZN(_13031_));
 AND2_X1 _22723_ (.A1(_11321_),
    .A2(_11427_),
    .ZN(_13032_));
 AOI211_X1 _22724_ (.A(_13031_),
    .B(_13032_),
    .C1(_11398_),
    .C2(_11427_),
    .ZN(_13033_));
 NAND2_X1 _22725_ (.A1(_11340_),
    .A2(_11414_),
    .ZN(_13034_));
 NAND2_X1 _22726_ (.A1(_13034_),
    .A2(_12308_),
    .ZN(_13035_));
 INV_X1 _22727_ (.A(_11361_),
    .ZN(_13036_));
 AND3_X1 _22728_ (.A1(_11380_),
    .A2(_13036_),
    .A3(_11414_),
    .ZN(_13037_));
 AOI211_X1 _22729_ (.A(_13035_),
    .B(_13037_),
    .C1(_11493_),
    .C2(_11414_),
    .ZN(_13038_));
 OAI21_X1 _22730_ (.A(_11431_),
    .B1(_11371_),
    .B2(_11525_),
    .ZN(_13039_));
 OAI211_X1 _22731_ (.A(_11427_),
    .B(_11373_),
    .C1(_11435_),
    .C2(_11335_),
    .ZN(_13040_));
 AND4_X1 _22732_ (.A1(_13033_),
    .A2(_13038_),
    .A3(_13039_),
    .A4(_13040_),
    .ZN(_13041_));
 NAND2_X1 _22733_ (.A1(_11409_),
    .A2(_11352_),
    .ZN(_13042_));
 NAND4_X1 _22734_ (.A1(_12670_),
    .A2(_12692_),
    .A3(_13042_),
    .A4(_11399_),
    .ZN(_13043_));
 AND2_X1 _22735_ (.A1(_11522_),
    .A2(_11423_),
    .ZN(_13044_));
 AND2_X1 _22736_ (.A1(_12717_),
    .A2(_11522_),
    .ZN(_13045_));
 OAI21_X1 _22737_ (.A(_12653_),
    .B1(_11523_),
    .B2(_12288_),
    .ZN(_13046_));
 NOR4_X1 _22738_ (.A1(_13043_),
    .A2(_13044_),
    .A3(_13045_),
    .A4(_13046_),
    .ZN(_13047_));
 AND2_X1 _22739_ (.A1(_11477_),
    .A2(_11467_),
    .ZN(_13048_));
 NOR2_X1 _22740_ (.A1(_11478_),
    .A2(_13048_),
    .ZN(_13049_));
 NAND2_X1 _22741_ (.A1(_12366_),
    .A2(_11370_),
    .ZN(_13050_));
 NAND4_X1 _22742_ (.A1(_13049_),
    .A2(_13050_),
    .A3(_12372_),
    .A4(_12668_),
    .ZN(_13051_));
 OAI211_X1 _22743_ (.A(_11382_),
    .B(_11396_),
    .C1(_11338_),
    .C2(_11360_),
    .ZN(_13052_));
 INV_X1 _22744_ (.A(_11382_),
    .ZN(_13053_));
 OAI21_X1 _22745_ (.A(_13052_),
    .B1(_12305_),
    .B2(_13053_),
    .ZN(_13054_));
 INV_X1 _22746_ (.A(_11418_),
    .ZN(_13055_));
 AND3_X1 _22747_ (.A1(_11363_),
    .A2(_11382_),
    .A3(_13055_),
    .ZN(_13056_));
 NAND2_X1 _22748_ (.A1(_11382_),
    .A2(_11429_),
    .ZN(_13057_));
 OAI21_X1 _22749_ (.A(_13057_),
    .B1(_13053_),
    .B2(_11526_),
    .ZN(_13058_));
 NOR4_X1 _22750_ (.A1(_13051_),
    .A2(_13054_),
    .A3(_13056_),
    .A4(_13058_),
    .ZN(_13059_));
 NAND4_X1 _22751_ (.A1(_13030_),
    .A2(_13041_),
    .A3(_13047_),
    .A4(_13059_),
    .ZN(_13060_));
 NAND2_X1 _22752_ (.A1(_11536_),
    .A2(_11437_),
    .ZN(_13061_));
 AOI21_X1 _22753_ (.A(_12313_),
    .B1(_11538_),
    .B2(_11539_),
    .ZN(_13062_));
 NAND2_X1 _22754_ (.A1(_11424_),
    .A2(_11487_),
    .ZN(_13063_));
 OAI211_X1 _22755_ (.A(_12315_),
    .B(_13063_),
    .C1(_12346_),
    .C2(_12313_),
    .ZN(_13064_));
 AOI211_X1 _22756_ (.A(_13062_),
    .B(_13064_),
    .C1(_11530_),
    .C2(_11488_),
    .ZN(_13065_));
 AND4_X1 _22757_ (.A1(_11389_),
    .A2(_11316_),
    .A3(_11343_),
    .A4(_11385_),
    .ZN(_13066_));
 NOR2_X1 _22758_ (.A1(_11535_),
    .A2(_13066_),
    .ZN(_13067_));
 OAI21_X1 _22759_ (.A(_11534_),
    .B1(_11346_),
    .B2(_11425_),
    .ZN(_13068_));
 AND4_X1 _22760_ (.A1(_13061_),
    .A2(_13065_),
    .A3(_13067_),
    .A4(_13068_),
    .ZN(_13069_));
 AND2_X1 _22761_ (.A1(_11334_),
    .A2(_11360_),
    .ZN(_13070_));
 OAI21_X1 _22762_ (.A(_11406_),
    .B1(_12375_),
    .B2(_13070_),
    .ZN(_13071_));
 AND2_X1 _22763_ (.A1(_11330_),
    .A2(_11473_),
    .ZN(_13072_));
 AOI211_X1 _22764_ (.A(_13072_),
    .B(_12681_),
    .C1(_11336_),
    .C2(_11331_),
    .ZN(_13073_));
 OAI21_X1 _22765_ (.A(_11406_),
    .B1(_11540_),
    .B2(_11321_),
    .ZN(_13074_));
 OAI21_X1 _22766_ (.A(_11347_),
    .B1(_12343_),
    .B2(_11400_),
    .ZN(_13075_));
 AND4_X1 _22767_ (.A1(_13071_),
    .A2(_13073_),
    .A3(_13074_),
    .A4(_13075_),
    .ZN(_13076_));
 OAI21_X1 _22768_ (.A(_11318_),
    .B1(_11452_),
    .B2(_11369_),
    .ZN(_13077_));
 OAI21_X1 _22769_ (.A(_13077_),
    .B1(_12318_),
    .B2(_11324_),
    .ZN(_13078_));
 AOI21_X1 _22770_ (.A(_11324_),
    .B1(_11441_),
    .B2(_12288_),
    .ZN(_13079_));
 AND2_X1 _22771_ (.A1(_12337_),
    .A2(_11318_),
    .ZN(_13080_));
 AND2_X1 _22772_ (.A1(_11318_),
    .A2(_12321_),
    .ZN(_13081_));
 NOR4_X1 _22773_ (.A1(_13078_),
    .A2(_13079_),
    .A3(_13080_),
    .A4(_13081_),
    .ZN(_13082_));
 OAI211_X1 _22774_ (.A(_11450_),
    .B(_11389_),
    .C1(_11338_),
    .C2(_11472_),
    .ZN(_13083_));
 AND2_X1 _22775_ (.A1(_11423_),
    .A2(_11360_),
    .ZN(_13084_));
 OAI21_X1 _22776_ (.A(_11450_),
    .B1(_11489_),
    .B2(_13084_),
    .ZN(_13085_));
 AND4_X1 _22777_ (.A1(_12336_),
    .A2(_13082_),
    .A3(_13083_),
    .A4(_13085_),
    .ZN(_13086_));
 AND2_X1 _22778_ (.A1(_11480_),
    .A2(_11429_),
    .ZN(_13087_));
 INV_X1 _22779_ (.A(_13087_),
    .ZN(_13088_));
 OAI21_X1 _22780_ (.A(_11481_),
    .B1(_11493_),
    .B2(_11528_),
    .ZN(_13089_));
 NAND3_X1 _22781_ (.A1(_11380_),
    .A2(_13036_),
    .A3(_11386_),
    .ZN(_13090_));
 NAND2_X1 _22782_ (.A1(_11425_),
    .A2(_11386_),
    .ZN(_13091_));
 AND4_X1 _22783_ (.A1(_13088_),
    .A2(_13089_),
    .A3(_13090_),
    .A4(_13091_),
    .ZN(_13092_));
 NAND4_X1 _22784_ (.A1(_13069_),
    .A2(_13076_),
    .A3(_13086_),
    .A4(_13092_),
    .ZN(_13093_));
 NOR2_X2 _22785_ (.A1(_13060_),
    .A2(_13093_),
    .ZN(_13094_));
 INV_X1 _22786_ (.A(_13094_),
    .ZN(_13095_));
 XNOR2_X1 _22787_ (.A(_13020_),
    .B(_13095_),
    .ZN(_13096_));
 XNOR2_X1 _22788_ (.A(_13019_),
    .B(_13096_),
    .ZN(_13097_));
 XNOR2_X1 _22789_ (.A(_13097_),
    .B(_17188_),
    .ZN(_13098_));
 MUX2_X1 _22790_ (.A(_12811_),
    .B(_13098_),
    .S(_11084_),
    .Z(_00719_));
 XOR2_X1 _22791_ (.A(_17189_),
    .B(_16992_),
    .Z(_13099_));
 AND4_X1 _22792_ (.A1(_11707_),
    .A2(_11732_),
    .A3(_11705_),
    .A4(_11588_),
    .ZN(_13100_));
 AND2_X1 _22793_ (.A1(_11777_),
    .A2(_11767_),
    .ZN(_13101_));
 AOI211_X1 _22794_ (.A(_13100_),
    .B(_13101_),
    .C1(_11644_),
    .C2(_11767_),
    .ZN(_13102_));
 OAI21_X1 _22795_ (.A(_11756_),
    .B1(_11598_),
    .B2(_12150_),
    .ZN(_13103_));
 OAI21_X1 _22796_ (.A(_11756_),
    .B1(_11737_),
    .B2(_11762_),
    .ZN(_13104_));
 AND4_X1 _22797_ (.A1(_11766_),
    .A2(_13102_),
    .A3(_13103_),
    .A4(_13104_),
    .ZN(_13105_));
 OAI21_X1 _22798_ (.A(_11675_),
    .B1(_11749_),
    .B2(_11694_),
    .ZN(_13106_));
 OAI211_X1 _22799_ (.A(_11675_),
    .B(_11709_),
    .C1(_11701_),
    .C2(_11661_),
    .ZN(_13107_));
 NAND2_X1 _22800_ (.A1(_12506_),
    .A2(_11675_),
    .ZN(_13108_));
 AND3_X1 _22801_ (.A1(_13106_),
    .A2(_13107_),
    .A3(_13108_),
    .ZN(_13109_));
 AND4_X1 _22802_ (.A1(_11642_),
    .A2(_11602_),
    .A3(_11571_),
    .A4(_11646_),
    .ZN(_13110_));
 NOR2_X1 _22803_ (.A1(_12522_),
    .A2(_11783_),
    .ZN(_13111_));
 AOI211_X1 _22804_ (.A(_13110_),
    .B(_13111_),
    .C1(_11639_),
    .C2(_11787_),
    .ZN(_13112_));
 OAI21_X1 _22805_ (.A(_11656_),
    .B1(_11768_),
    .B2(_11657_),
    .ZN(_13113_));
 AND3_X1 _22806_ (.A1(_13113_),
    .A2(_11651_),
    .A3(_12168_),
    .ZN(_13114_));
 AND2_X1 _22807_ (.A1(_11821_),
    .A2(_11694_),
    .ZN(_13115_));
 NOR4_X1 _22808_ (.A1(_11663_),
    .A2(_12165_),
    .A3(_12888_),
    .A4(_13115_),
    .ZN(_13116_));
 AND4_X1 _22809_ (.A1(_13109_),
    .A2(_13112_),
    .A3(_13114_),
    .A4(_13116_),
    .ZN(_13117_));
 AND4_X1 _22810_ (.A1(_11824_),
    .A2(_11702_),
    .A3(_11732_),
    .A4(_11572_),
    .ZN(_13118_));
 AOI211_X1 _22811_ (.A(_13118_),
    .B(_12563_),
    .C1(_11577_),
    .C2(_12122_),
    .ZN(_13119_));
 INV_X1 _22812_ (.A(_11792_),
    .ZN(_13120_));
 INV_X1 _22813_ (.A(_11791_),
    .ZN(_13121_));
 NAND2_X1 _22814_ (.A1(_11735_),
    .A2(_11577_),
    .ZN(_13122_));
 OAI21_X1 _22815_ (.A(_11735_),
    .B1(_11725_),
    .B2(_11644_),
    .ZN(_13123_));
 AND4_X1 _22816_ (.A1(_13120_),
    .A2(_13121_),
    .A3(_13122_),
    .A4(_13123_),
    .ZN(_13124_));
 AND4_X1 _22817_ (.A1(_13105_),
    .A2(_13117_),
    .A3(_13119_),
    .A4(_13124_),
    .ZN(_13125_));
 AND2_X1 _22818_ (.A1(_11581_),
    .A2(_11604_),
    .ZN(_13126_));
 INV_X1 _22819_ (.A(_13126_),
    .ZN(_13127_));
 OAI211_X1 _22820_ (.A(_13127_),
    .B(_11835_),
    .C1(_11591_),
    .C2(_11758_),
    .ZN(_13128_));
 OR2_X1 _22821_ (.A1(_11829_),
    .A2(_11830_),
    .ZN(_13129_));
 AOI21_X1 _22822_ (.A(_11591_),
    .B1(_11746_),
    .B2(_11840_),
    .ZN(_13130_));
 OAI211_X1 _22823_ (.A(_11566_),
    .B(_11659_),
    .C1(_11563_),
    .C2(_11564_),
    .ZN(_13131_));
 NAND2_X1 _22824_ (.A1(_12149_),
    .A2(_11683_),
    .ZN(_13132_));
 NAND4_X1 _22825_ (.A1(_11669_),
    .A2(_11671_),
    .A3(_11566_),
    .A4(_11659_),
    .ZN(_13133_));
 NAND4_X1 _22826_ (.A1(_13131_),
    .A2(_12942_),
    .A3(_13132_),
    .A4(_13133_),
    .ZN(_13134_));
 NOR4_X1 _22827_ (.A1(_13128_),
    .A2(_13129_),
    .A3(_13130_),
    .A4(_13134_),
    .ZN(_13135_));
 NAND2_X1 _22828_ (.A1(_11680_),
    .A2(_11612_),
    .ZN(_13136_));
 AOI211_X1 _22829_ (.A(_12929_),
    .B(_12133_),
    .C1(_11777_),
    .C2(_11680_),
    .ZN(_13137_));
 NAND2_X1 _22830_ (.A1(_12150_),
    .A2(_11714_),
    .ZN(_13138_));
 NAND3_X1 _22831_ (.A1(_11714_),
    .A2(_11702_),
    .A3(_11710_),
    .ZN(_13139_));
 NAND2_X1 _22832_ (.A1(_11689_),
    .A2(_11714_),
    .ZN(_13140_));
 AND4_X1 _22833_ (.A1(_13138_),
    .A2(_12524_),
    .A3(_13139_),
    .A4(_13140_),
    .ZN(_13141_));
 OAI211_X1 _22834_ (.A(_11680_),
    .B(_11702_),
    .C1(_11706_),
    .C2(_11707_),
    .ZN(_13142_));
 AND4_X1 _22835_ (.A1(_13136_),
    .A2(_13137_),
    .A3(_13141_),
    .A4(_13142_),
    .ZN(_13143_));
 OAI211_X1 _22836_ (.A(_11606_),
    .B(_11611_),
    .C1(_11682_),
    .C2(_11843_),
    .ZN(_13144_));
 NAND2_X1 _22837_ (.A1(_11553_),
    .A2(_11557_),
    .ZN(_13145_));
 NAND4_X1 _22838_ (.A1(_11566_),
    .A2(_11592_),
    .A3(_11583_),
    .A4(_11572_),
    .ZN(_13146_));
 OAI211_X1 _22839_ (.A(_13145_),
    .B(_13146_),
    .C1(_11847_),
    .C2(_11684_),
    .ZN(_13147_));
 AOI21_X1 _22840_ (.A(_11843_),
    .B1(_11860_),
    .B2(_11741_),
    .ZN(_13148_));
 NOR4_X1 _22841_ (.A1(_13144_),
    .A2(_12147_),
    .A3(_13147_),
    .A4(_13148_),
    .ZN(_13149_));
 OAI21_X1 _22842_ (.A(_11722_),
    .B1(_11689_),
    .B2(_11587_),
    .ZN(_13150_));
 OAI211_X1 _22843_ (.A(_11704_),
    .B(_11702_),
    .C1(_11706_),
    .C2(_11707_),
    .ZN(_13151_));
 NAND2_X1 _22844_ (.A1(_11704_),
    .A2(_11644_),
    .ZN(_13152_));
 NAND4_X1 _22845_ (.A1(_11709_),
    .A2(_11661_),
    .A3(_11695_),
    .A4(_11588_),
    .ZN(_13153_));
 AND3_X1 _22846_ (.A1(_13151_),
    .A2(_13152_),
    .A3(_13153_),
    .ZN(_13154_));
 OAI21_X1 _22847_ (.A(_11722_),
    .B1(_11720_),
    .B2(_11640_),
    .ZN(_13155_));
 OAI211_X1 _22848_ (.A(_11695_),
    .B(_11659_),
    .C1(_11564_),
    .C2(_11644_),
    .ZN(_13156_));
 AND4_X1 _22849_ (.A1(_13150_),
    .A2(_13154_),
    .A3(_13155_),
    .A4(_13156_),
    .ZN(_13157_));
 AND4_X1 _22850_ (.A1(_13135_),
    .A2(_13143_),
    .A3(_13149_),
    .A4(_13157_),
    .ZN(_13158_));
 AND2_X1 _22851_ (.A1(_13125_),
    .A2(_13158_),
    .ZN(_13159_));
 AND2_X1 _22852_ (.A1(_12264_),
    .A2(_11270_),
    .ZN(_13160_));
 AOI21_X1 _22853_ (.A(_12266_),
    .B1(_11277_),
    .B2(_12260_),
    .ZN(_13161_));
 AND4_X1 _22854_ (.A1(_11150_),
    .A2(_11238_),
    .A3(_11141_),
    .A4(_12182_),
    .ZN(_13162_));
 NOR3_X1 _22855_ (.A1(_13160_),
    .A2(_13161_),
    .A3(_13162_),
    .ZN(_13163_));
 NAND4_X1 _22856_ (.A1(_13163_),
    .A2(_11236_),
    .A3(_12270_),
    .A4(_12610_),
    .ZN(_13164_));
 OAI21_X1 _22857_ (.A(_11285_),
    .B1(_11181_),
    .B2(_11132_),
    .ZN(_13165_));
 OAI21_X1 _22858_ (.A(_11285_),
    .B1(_11302_),
    .B2(_11286_),
    .ZN(_13166_));
 OAI21_X1 _22859_ (.A(_11299_),
    .B1(_12829_),
    .B2(_11185_),
    .ZN(_13167_));
 NAND4_X1 _22860_ (.A1(_13165_),
    .A2(_13166_),
    .A3(_13167_),
    .A4(_11298_),
    .ZN(_13168_));
 OAI21_X1 _22861_ (.A(_11247_),
    .B1(_11269_),
    .B2(_12580_),
    .ZN(_13169_));
 OAI21_X1 _22862_ (.A(_11259_),
    .B1(_11267_),
    .B2(_12275_),
    .ZN(_13170_));
 AND2_X1 _22863_ (.A1(_13170_),
    .A2(_12877_),
    .ZN(_13171_));
 NAND4_X1 _22864_ (.A1(_13169_),
    .A2(_11257_),
    .A3(_11256_),
    .A4(_13171_),
    .ZN(_13172_));
 NAND2_X1 _22865_ (.A1(_11267_),
    .A2(_11264_),
    .ZN(_13173_));
 NAND2_X1 _22866_ (.A1(_12205_),
    .A2(_11264_),
    .ZN(_13174_));
 NAND2_X1 _22867_ (.A1(_13173_),
    .A2(_13174_),
    .ZN(_13175_));
 AND2_X1 _22868_ (.A1(_11264_),
    .A2(_11160_),
    .ZN(_13176_));
 NOR2_X1 _22869_ (.A1(_13175_),
    .A2(_13176_),
    .ZN(_13177_));
 OAI21_X1 _22870_ (.A(_11295_),
    .B1(_12221_),
    .B2(_11160_),
    .ZN(_13178_));
 OAI21_X1 _22871_ (.A(_11265_),
    .B1(_11225_),
    .B2(_11235_),
    .ZN(_13179_));
 NAND4_X1 _22872_ (.A1(_13177_),
    .A2(_12586_),
    .A3(_13178_),
    .A4(_13179_),
    .ZN(_13180_));
 NOR4_X1 _22873_ (.A1(_13164_),
    .A2(_13168_),
    .A3(_13172_),
    .A4(_13180_),
    .ZN(_13181_));
 OAI21_X1 _22874_ (.A(_11093_),
    .B1(_11279_),
    .B2(_12205_),
    .ZN(_13182_));
 NAND2_X1 _22875_ (.A1(_11093_),
    .A2(_11162_),
    .ZN(_13183_));
 OAI21_X1 _22876_ (.A(_11093_),
    .B1(_11121_),
    .B2(_11139_),
    .ZN(_13184_));
 NAND3_X1 _22877_ (.A1(_13182_),
    .A2(_13183_),
    .A3(_13184_),
    .ZN(_13185_));
 AND2_X1 _22878_ (.A1(_11301_),
    .A2(_11103_),
    .ZN(_13186_));
 AND2_X1 _22879_ (.A1(_11103_),
    .A2(_12187_),
    .ZN(_13187_));
 NOR2_X1 _22880_ (.A1(_13186_),
    .A2(_13187_),
    .ZN(_13188_));
 INV_X1 _22881_ (.A(_13188_),
    .ZN(_13189_));
 AOI21_X1 _22882_ (.A(_11107_),
    .B1(_11293_),
    .B2(_11218_),
    .ZN(_13190_));
 NAND2_X1 _22883_ (.A1(_11152_),
    .A2(_11129_),
    .ZN(_13191_));
 NAND4_X1 _22884_ (.A1(_11091_),
    .A2(_11189_),
    .A3(_11195_),
    .A4(_11239_),
    .ZN(_13192_));
 OAI211_X1 _22885_ (.A(_13191_),
    .B(_13192_),
    .C1(_11283_),
    .C2(_11107_),
    .ZN(_13193_));
 NOR4_X1 _22886_ (.A1(_13185_),
    .A2(_13189_),
    .A3(_13190_),
    .A4(_13193_),
    .ZN(_13194_));
 OAI21_X1 _22887_ (.A(_11221_),
    .B1(_11204_),
    .B2(_11185_),
    .ZN(_13195_));
 OAI211_X1 _22888_ (.A(_11199_),
    .B(_11100_),
    .C1(_11109_),
    .C2(_11142_),
    .ZN(_13196_));
 OAI21_X1 _22889_ (.A(_11199_),
    .B1(_12829_),
    .B2(_11235_),
    .ZN(_13197_));
 OAI21_X1 _22890_ (.A(_11221_),
    .B1(_11220_),
    .B2(_11223_),
    .ZN(_13198_));
 AND4_X1 _22891_ (.A1(_13195_),
    .A2(_13196_),
    .A3(_13197_),
    .A4(_13198_),
    .ZN(_13199_));
 OAI211_X1 _22892_ (.A(_11137_),
    .B(_11100_),
    .C1(_11189_),
    .C2(_11155_),
    .ZN(_13200_));
 NAND4_X1 _22893_ (.A1(_11091_),
    .A2(_11115_),
    .A3(_11143_),
    .A4(_11239_),
    .ZN(_13201_));
 NAND3_X1 _22894_ (.A1(_12213_),
    .A2(_13200_),
    .A3(_13201_),
    .ZN(_13202_));
 AOI21_X1 _22895_ (.A(_12224_),
    .B1(_12589_),
    .B2(_11178_),
    .ZN(_13203_));
 OAI21_X1 _22896_ (.A(_12834_),
    .B1(_12224_),
    .B2(_11122_),
    .ZN(_13204_));
 AND2_X1 _22897_ (.A1(_11149_),
    .A2(_11160_),
    .ZN(_13205_));
 NOR4_X1 _22898_ (.A1(_13202_),
    .A2(_13203_),
    .A3(_13204_),
    .A4(_13205_),
    .ZN(_13206_));
 OAI21_X1 _22899_ (.A(_11175_),
    .B1(_11159_),
    .B2(_11190_),
    .ZN(_13207_));
 NAND2_X1 _22900_ (.A1(_12829_),
    .A2(_11207_),
    .ZN(_13208_));
 AND3_X1 _22901_ (.A1(_12243_),
    .A2(_13208_),
    .A3(_12816_),
    .ZN(_13209_));
 NAND2_X1 _22902_ (.A1(_11207_),
    .A2(_11105_),
    .ZN(_13210_));
 NAND4_X1 _22903_ (.A1(_11194_),
    .A2(_12182_),
    .A3(_11115_),
    .A4(_11193_),
    .ZN(_13211_));
 AND3_X1 _22904_ (.A1(_12814_),
    .A2(_13210_),
    .A3(_13211_),
    .ZN(_13212_));
 OAI21_X1 _22905_ (.A(_11175_),
    .B1(_12199_),
    .B2(_12642_),
    .ZN(_13213_));
 AND4_X1 _22906_ (.A1(_13207_),
    .A2(_13209_),
    .A3(_13212_),
    .A4(_13213_),
    .ZN(_13214_));
 AND4_X1 _22907_ (.A1(_13194_),
    .A2(_13199_),
    .A3(_13206_),
    .A4(_13214_),
    .ZN(_13215_));
 AND2_X2 _22908_ (.A1(_13181_),
    .A2(_13215_),
    .ZN(_13216_));
 XOR2_X2 _22909_ (.A(_13159_),
    .B(_13216_),
    .Z(_13217_));
 OAI21_X1 _22910_ (.A(_12480_),
    .B1(_12041_),
    .B2(_12080_),
    .ZN(_13218_));
 NAND2_X1 _22911_ (.A1(_12480_),
    .A2(_12412_),
    .ZN(_13219_));
 AND3_X1 _22912_ (.A1(_13218_),
    .A2(_11965_),
    .A3(_13219_),
    .ZN(_13220_));
 NAND3_X1 _22913_ (.A1(_11943_),
    .A2(_11906_),
    .A3(_11944_),
    .ZN(_13221_));
 NAND2_X1 _22914_ (.A1(_12447_),
    .A2(_11943_),
    .ZN(_13222_));
 OAI211_X1 _22915_ (.A(_13221_),
    .B(_13222_),
    .C1(_12432_),
    .C2(_12753_),
    .ZN(_13223_));
 AOI21_X1 _22916_ (.A(_12753_),
    .B1(_12387_),
    .B2(_12999_),
    .ZN(_13224_));
 NOR4_X1 _22917_ (.A1(_13223_),
    .A2(_13224_),
    .A3(_12473_),
    .A4(_11949_),
    .ZN(_13225_));
 OAI211_X1 _22918_ (.A(_12489_),
    .B(_12414_),
    .C1(_11919_),
    .C2(_11906_),
    .ZN(_13226_));
 OAI211_X1 _22919_ (.A(_12489_),
    .B(_12010_),
    .C1(_11945_),
    .C2(_11946_),
    .ZN(_13227_));
 OAI21_X1 _22920_ (.A(_12489_),
    .B1(_11987_),
    .B2(_12401_),
    .ZN(_13228_));
 AND4_X1 _22921_ (.A1(_12490_),
    .A2(_13226_),
    .A3(_13227_),
    .A4(_13228_),
    .ZN(_13229_));
 OAI211_X1 _22922_ (.A(_12762_),
    .B(_11955_),
    .C1(_11927_),
    .C2(_11920_),
    .ZN(_13230_));
 OAI211_X1 _22923_ (.A(_12762_),
    .B(_12414_),
    .C1(_11932_),
    .C2(_11933_),
    .ZN(_13231_));
 OAI211_X1 _22924_ (.A(_12762_),
    .B(_12010_),
    .C1(_11945_),
    .C2(_11933_),
    .ZN(_13232_));
 OAI21_X1 _22925_ (.A(_12762_),
    .B1(_12410_),
    .B2(_12412_),
    .ZN(_13233_));
 AND4_X1 _22926_ (.A1(_13230_),
    .A2(_13231_),
    .A3(_13232_),
    .A4(_13233_),
    .ZN(_13234_));
 NAND4_X1 _22927_ (.A1(_13220_),
    .A2(_13225_),
    .A3(_13229_),
    .A4(_13234_),
    .ZN(_13235_));
 NAND2_X1 _22928_ (.A1(_12006_),
    .A2(_12033_),
    .ZN(_13236_));
 AND2_X1 _22929_ (.A1(_12467_),
    .A2(_13236_),
    .ZN(_13237_));
 INV_X1 _22930_ (.A(_13237_),
    .ZN(_13238_));
 AND2_X1 _22931_ (.A1(_12009_),
    .A2(_12763_),
    .ZN(_13239_));
 AND2_X1 _22932_ (.A1(_12009_),
    .A2(_11980_),
    .ZN(_13240_));
 NOR4_X1 _22933_ (.A1(_13238_),
    .A2(_13239_),
    .A3(_13240_),
    .A4(_12775_),
    .ZN(_13241_));
 AND4_X1 _22934_ (.A1(_11946_),
    .A2(_11978_),
    .A3(_11924_),
    .A4(_12011_),
    .ZN(_13242_));
 AND2_X1 _22935_ (.A1(_12461_),
    .A2(_11953_),
    .ZN(_13243_));
 AOI211_X1 _22936_ (.A(_13242_),
    .B(_13243_),
    .C1(_12461_),
    .C2(_12389_),
    .ZN(_13244_));
 NAND4_X1 _22937_ (.A1(_11979_),
    .A2(_11945_),
    .A3(_11955_),
    .A4(_11924_),
    .ZN(_13245_));
 OAI211_X1 _22938_ (.A(_12461_),
    .B(_12414_),
    .C1(_11932_),
    .C2(_11946_),
    .ZN(_13246_));
 NAND4_X1 _22939_ (.A1(_13241_),
    .A2(_13244_),
    .A3(_13245_),
    .A4(_13246_),
    .ZN(_13247_));
 AND2_X1 _22940_ (.A1(_12394_),
    .A2(_11993_),
    .ZN(_13248_));
 AND2_X1 _22941_ (.A1(_11993_),
    .A2(_12034_),
    .ZN(_13249_));
 AND2_X1 _22942_ (.A1(_11993_),
    .A2(_12001_),
    .ZN(_13250_));
 OR4_X1 _22943_ (.A1(_12963_),
    .A2(_13248_),
    .A3(_13249_),
    .A4(_13250_),
    .ZN(_13251_));
 AND3_X1 _22944_ (.A1(_12449_),
    .A2(_11957_),
    .A3(_11978_),
    .ZN(_13252_));
 OR4_X1 _22945_ (.A1(_11975_),
    .A2(_12801_),
    .A3(_12960_),
    .A4(_13252_),
    .ZN(_13253_));
 NOR4_X1 _22946_ (.A1(_13235_),
    .A2(_13247_),
    .A3(_13251_),
    .A4(_13253_),
    .ZN(_13254_));
 AOI21_X1 _22947_ (.A(_12037_),
    .B1(_12400_),
    .B2(_12075_),
    .ZN(_13255_));
 AND3_X1 _22948_ (.A1(_12391_),
    .A2(_12010_),
    .A3(_11919_),
    .ZN(_13256_));
 AND2_X1 _22949_ (.A1(_12410_),
    .A2(_12391_),
    .ZN(_13257_));
 NOR4_X1 _22950_ (.A1(_13255_),
    .A2(_12031_),
    .A3(_13256_),
    .A4(_13257_),
    .ZN(_13258_));
 NOR2_X1 _22951_ (.A1(_12044_),
    .A2(_12459_),
    .ZN(_13259_));
 AOI21_X1 _22952_ (.A(_13259_),
    .B1(_11937_),
    .B2(_12022_),
    .ZN(_13260_));
 AND3_X1 _22953_ (.A1(_12410_),
    .A2(_12018_),
    .A3(_11977_),
    .ZN(_13261_));
 AOI21_X1 _22954_ (.A(_13261_),
    .B1(_12389_),
    .B2(_12022_),
    .ZN(_13262_));
 NAND2_X1 _22955_ (.A1(_11953_),
    .A2(_12094_),
    .ZN(_13263_));
 OAI21_X1 _22956_ (.A(_12089_),
    .B1(_12033_),
    .B2(_12034_),
    .ZN(_13264_));
 OAI21_X1 _22957_ (.A(_12094_),
    .B1(_12080_),
    .B2(_12449_),
    .ZN(_13265_));
 NAND2_X1 _22958_ (.A1(_11907_),
    .A2(_12088_),
    .ZN(_13266_));
 AND4_X1 _22959_ (.A1(_13263_),
    .A2(_13264_),
    .A3(_13265_),
    .A4(_13266_),
    .ZN(_13267_));
 NAND4_X1 _22960_ (.A1(_13258_),
    .A2(_13260_),
    .A3(_13262_),
    .A4(_13267_),
    .ZN(_13268_));
 OAI21_X1 _22961_ (.A(_12440_),
    .B1(_12399_),
    .B2(_12447_),
    .ZN(_13269_));
 AND2_X1 _22962_ (.A1(_11918_),
    .A2(_11932_),
    .ZN(_13270_));
 INV_X1 _22963_ (.A(_13270_),
    .ZN(_13271_));
 OAI211_X1 _22964_ (.A(_13269_),
    .B(_12990_),
    .C1(_12445_),
    .C2(_13271_),
    .ZN(_13272_));
 NAND2_X1 _22965_ (.A1(_12064_),
    .A2(_12425_),
    .ZN(_13273_));
 NAND2_X1 _22966_ (.A1(_11898_),
    .A2(_12423_),
    .ZN(_13274_));
 OAI21_X1 _22967_ (.A(_12064_),
    .B1(_11953_),
    .B2(_12412_),
    .ZN(_13275_));
 NAND4_X1 _22968_ (.A1(_12795_),
    .A2(_13273_),
    .A3(_13274_),
    .A4(_13275_),
    .ZN(_13276_));
 OR2_X1 _22969_ (.A1(_13272_),
    .A2(_13276_),
    .ZN(_13277_));
 OAI211_X1 _22970_ (.A(_12078_),
    .B(_11955_),
    .C1(_11932_),
    .C2(_11946_),
    .ZN(_13278_));
 OAI21_X1 _22971_ (.A(_12078_),
    .B1(_11929_),
    .B2(_11930_),
    .ZN(_13279_));
 OAI211_X1 _22972_ (.A(_13278_),
    .B(_13279_),
    .C1(_12079_),
    .C2(_12398_),
    .ZN(_13280_));
 AND2_X1 _22973_ (.A1(_12068_),
    .A2(_12449_),
    .ZN(_13281_));
 AOI21_X1 _22974_ (.A(_12069_),
    .B1(_12083_),
    .B2(_12999_),
    .ZN(_13282_));
 AND2_X1 _22975_ (.A1(_12068_),
    .A2(_11985_),
    .ZN(_13283_));
 AND3_X1 _22976_ (.A1(_11957_),
    .A2(_12049_),
    .A3(_12011_),
    .ZN(_13284_));
 OR4_X1 _22977_ (.A1(_13281_),
    .A2(_13282_),
    .A3(_13283_),
    .A4(_13284_),
    .ZN(_13285_));
 NOR4_X1 _22978_ (.A1(_13268_),
    .A2(_13277_),
    .A3(_13280_),
    .A4(_13285_),
    .ZN(_13286_));
 AND2_X2 _22979_ (.A1(_13254_),
    .A2(_13286_),
    .ZN(_13287_));
 XNOR2_X1 _22980_ (.A(_13287_),
    .B(_12102_),
    .ZN(_13288_));
 XNOR2_X1 _22981_ (.A(_13217_),
    .B(_13288_),
    .ZN(_13289_));
 XOR2_X2 _22982_ (.A(_11877_),
    .B(_12952_),
    .Z(_13290_));
 OAI211_X1 _22983_ (.A(_11347_),
    .B(_11423_),
    .C1(_11435_),
    .C2(_11472_),
    .ZN(_13291_));
 NAND3_X1 _22984_ (.A1(_11347_),
    .A2(_13036_),
    .A3(_12690_),
    .ZN(_13292_));
 NAND4_X1 _22985_ (.A1(_13291_),
    .A2(_11337_),
    .A3(_11500_),
    .A4(_13292_),
    .ZN(_13293_));
 AOI21_X1 _22986_ (.A(_12697_),
    .B1(_12318_),
    .B2(_11526_),
    .ZN(_13294_));
 AOI21_X1 _22987_ (.A(_12697_),
    .B1(_11378_),
    .B2(_11443_),
    .ZN(_13295_));
 AND3_X1 _22988_ (.A1(_11405_),
    .A2(_11408_),
    .A3(_11334_),
    .ZN(_13296_));
 NOR4_X1 _22989_ (.A1(_13293_),
    .A2(_13294_),
    .A3(_13295_),
    .A4(_13296_),
    .ZN(_13297_));
 OAI21_X1 _22990_ (.A(_11482_),
    .B1(_11410_),
    .B2(_11344_),
    .ZN(_13298_));
 AND3_X1 _22991_ (.A1(_11483_),
    .A2(_11362_),
    .A3(_11373_),
    .ZN(_13299_));
 AOI21_X1 _22992_ (.A(_11387_),
    .B1(_12346_),
    .B2(_12724_),
    .ZN(_13300_));
 AOI211_X1 _22993_ (.A(_13299_),
    .B(_13300_),
    .C1(_11483_),
    .C2(_11380_),
    .ZN(_13301_));
 OAI221_X1 _22994_ (.A(_11482_),
    .B1(_11435_),
    .B2(_11418_),
    .C1(_11396_),
    .C2(_11389_),
    .ZN(_13302_));
 OAI211_X1 _22995_ (.A(_11385_),
    .B(_11364_),
    .C1(_11371_),
    .C2(_11525_),
    .ZN(_13303_));
 AND4_X1 _22996_ (.A1(_13298_),
    .A2(_13301_),
    .A3(_13302_),
    .A4(_13303_),
    .ZN(_13304_));
 INV_X1 _22997_ (.A(_11497_),
    .ZN(_13305_));
 OAI21_X1 _22998_ (.A(_11498_),
    .B1(_11538_),
    .B2(_13305_),
    .ZN(_13306_));
 AOI21_X1 _22999_ (.A(_13306_),
    .B1(_11321_),
    .B2(_11497_),
    .ZN(_13307_));
 NAND2_X1 _23000_ (.A1(_11403_),
    .A2(_11327_),
    .ZN(_13308_));
 AND3_X1 _23001_ (.A1(_12671_),
    .A2(_11519_),
    .A3(_13308_),
    .ZN(_13309_));
 OAI21_X1 _23002_ (.A(_11403_),
    .B1(_11452_),
    .B2(_12322_),
    .ZN(_13310_));
 AND4_X1 _23003_ (.A1(_12339_),
    .A2(_13307_),
    .A3(_13309_),
    .A4(_13310_),
    .ZN(_13311_));
 NAND2_X1 _23004_ (.A1(_12343_),
    .A2(_11487_),
    .ZN(_13312_));
 NAND2_X1 _23005_ (.A1(_11534_),
    .A2(_11321_),
    .ZN(_13313_));
 OAI21_X1 _23006_ (.A(_11536_),
    .B1(_11452_),
    .B2(_11425_),
    .ZN(_13314_));
 NAND2_X1 _23007_ (.A1(_11380_),
    .A2(_11533_),
    .ZN(_13315_));
 NAND2_X1 _23008_ (.A1(_11489_),
    .A2(_11534_),
    .ZN(_13316_));
 AND4_X1 _23009_ (.A1(_13313_),
    .A2(_13314_),
    .A3(_13315_),
    .A4(_13316_),
    .ZN(_13317_));
 NAND3_X1 _23010_ (.A1(_11488_),
    .A2(_11396_),
    .A3(_11343_),
    .ZN(_13318_));
 OAI21_X1 _23011_ (.A(_11488_),
    .B1(_12664_),
    .B2(_11344_),
    .ZN(_13319_));
 AND4_X1 _23012_ (.A1(_13312_),
    .A2(_13317_),
    .A3(_13318_),
    .A4(_13319_),
    .ZN(_13320_));
 AND4_X1 _23013_ (.A1(_13297_),
    .A2(_13304_),
    .A3(_13311_),
    .A4(_13320_),
    .ZN(_13321_));
 OAI21_X1 _23014_ (.A(_11434_),
    .B1(_12343_),
    .B2(_11528_),
    .ZN(_13322_));
 OAI211_X1 _23015_ (.A(_11460_),
    .B(_16746_),
    .C1(_16745_),
    .C2(_11362_),
    .ZN(_13323_));
 OAI21_X1 _23016_ (.A(_11434_),
    .B1(_12338_),
    .B2(_11456_),
    .ZN(_13324_));
 AND4_X1 _23017_ (.A1(_11502_),
    .A2(_13322_),
    .A3(_13323_),
    .A4(_13324_),
    .ZN(_13325_));
 OAI21_X1 _23018_ (.A(_12374_),
    .B1(_12717_),
    .B2(_12375_),
    .ZN(_13326_));
 OAI21_X1 _23019_ (.A(_13326_),
    .B1(_11421_),
    .B2(_13053_),
    .ZN(_13327_));
 NAND3_X1 _23020_ (.A1(_11420_),
    .A2(_11364_),
    .A3(_11368_),
    .ZN(_13328_));
 NAND2_X1 _23021_ (.A1(_12371_),
    .A2(_13328_),
    .ZN(_13329_));
 NOR4_X1 _23022_ (.A1(_13327_),
    .A2(_11375_),
    .A3(_13329_),
    .A4(_13048_),
    .ZN(_13330_));
 AND2_X1 _23023_ (.A1(_11419_),
    .A2(_11414_),
    .ZN(_13331_));
 INV_X1 _23024_ (.A(_13331_),
    .ZN(_13332_));
 AND2_X1 _23025_ (.A1(_11499_),
    .A2(_11413_),
    .ZN(_13333_));
 INV_X1 _23026_ (.A(_13333_),
    .ZN(_13334_));
 NAND2_X1 _23027_ (.A1(_11415_),
    .A2(_11327_),
    .ZN(_13335_));
 AND3_X1 _23028_ (.A1(_13332_),
    .A2(_13334_),
    .A3(_13335_),
    .ZN(_13336_));
 AOI21_X1 _23029_ (.A(_13035_),
    .B1(_11415_),
    .B2(_12717_),
    .ZN(_13337_));
 OAI21_X1 _23030_ (.A(_11431_),
    .B1(_12324_),
    .B2(_11327_),
    .ZN(_13338_));
 AND4_X1 _23031_ (.A1(_12687_),
    .A2(_13336_),
    .A3(_13337_),
    .A4(_13338_),
    .ZN(_13339_));
 NAND2_X1 _23032_ (.A1(_13044_),
    .A2(_13055_),
    .ZN(_13340_));
 OAI21_X1 _23033_ (.A(_11522_),
    .B1(_11511_),
    .B2(_11321_),
    .ZN(_13341_));
 NAND4_X1 _23034_ (.A1(_11368_),
    .A2(_11316_),
    .A3(_11373_),
    .A4(_11338_),
    .ZN(_13342_));
 NAND3_X1 _23035_ (.A1(_13340_),
    .A2(_13341_),
    .A3(_13342_),
    .ZN(_13343_));
 NOR4_X1 _23036_ (.A1(_13343_),
    .A2(_12362_),
    .A3(_11357_),
    .A4(_12669_),
    .ZN(_13344_));
 AND4_X1 _23037_ (.A1(_13325_),
    .A2(_13330_),
    .A3(_13339_),
    .A4(_13344_),
    .ZN(_13345_));
 NAND2_X2 _23038_ (.A1(_13321_),
    .A2(_13345_),
    .ZN(_13346_));
 XNOR2_X1 _23039_ (.A(_13290_),
    .B(_13346_),
    .ZN(_13347_));
 XNOR2_X1 _23040_ (.A(_13289_),
    .B(_13347_),
    .ZN(_13348_));
 XNOR2_X1 _23041_ (.A(_13348_),
    .B(_17189_),
    .ZN(_13349_));
 MUX2_X1 _23042_ (.A(_13099_),
    .B(_13349_),
    .S(_11084_),
    .Z(_00720_));
 XOR2_X1 _23043_ (.A(_17190_),
    .B(_16993_),
    .Z(_13350_));
 OAI21_X1 _23044_ (.A(_11093_),
    .B1(_12205_),
    .B2(_11190_),
    .ZN(_13351_));
 AND2_X1 _23045_ (.A1(_11116_),
    .A2(_11103_),
    .ZN(_13352_));
 AOI211_X1 _23046_ (.A(_13352_),
    .B(_13186_),
    .C1(_12617_),
    .C2(_11129_),
    .ZN(_13353_));
 OAI21_X1 _23047_ (.A(_11093_),
    .B1(_11162_),
    .B2(_11286_),
    .ZN(_13354_));
 OAI21_X1 _23048_ (.A(_11129_),
    .B1(_12275_),
    .B2(_11152_),
    .ZN(_13355_));
 AND4_X1 _23049_ (.A1(_13351_),
    .A2(_13353_),
    .A3(_13354_),
    .A4(_13355_),
    .ZN(_13356_));
 OAI21_X1 _23050_ (.A(_11137_),
    .B1(_11267_),
    .B2(_11133_),
    .ZN(_13357_));
 OAI211_X1 _23051_ (.A(_11149_),
    .B(_11194_),
    .C1(_11109_),
    .C2(_11173_),
    .ZN(_13358_));
 OAI211_X1 _23052_ (.A(_11149_),
    .B(_11141_),
    .C1(_11150_),
    .C2(_11173_),
    .ZN(_13359_));
 AND3_X1 _23053_ (.A1(_13358_),
    .A2(_13359_),
    .A3(_12837_),
    .ZN(_13360_));
 AND4_X1 _23054_ (.A1(_11146_),
    .A2(_13356_),
    .A3(_13357_),
    .A4(_13360_),
    .ZN(_13361_));
 AOI21_X1 _23055_ (.A(_12250_),
    .B1(_11293_),
    .B2(_11218_),
    .ZN(_13362_));
 AND2_X1 _23056_ (.A1(_11116_),
    .A2(_11199_),
    .ZN(_13363_));
 AND4_X1 _23057_ (.A1(_11193_),
    .A2(_11155_),
    .A3(_11239_),
    .A4(_11195_),
    .ZN(_13364_));
 NOR3_X1 _23058_ (.A1(_13362_),
    .A2(_13363_),
    .A3(_13364_),
    .ZN(_13365_));
 AOI221_X1 _23059_ (.A(_11172_),
    .B1(_11109_),
    .B2(_11186_),
    .C1(_12198_),
    .C2(_11169_),
    .ZN(_13366_));
 AOI211_X1 _23060_ (.A(_12246_),
    .B(_13366_),
    .C1(_11175_),
    .C2(_11190_),
    .ZN(_13367_));
 OAI21_X1 _23061_ (.A(_11207_),
    .B1(_12617_),
    .B2(_11273_),
    .ZN(_13368_));
 NAND2_X1 _23062_ (.A1(_12864_),
    .A2(_11207_),
    .ZN(_13369_));
 AND3_X1 _23063_ (.A1(_13368_),
    .A2(_13210_),
    .A3(_13369_),
    .ZN(_13370_));
 AOI21_X1 _23064_ (.A(_11214_),
    .B1(_12251_),
    .B2(_12219_),
    .ZN(_13371_));
 AND2_X1 _23065_ (.A1(_11220_),
    .A2(_11221_),
    .ZN(_13372_));
 AND4_X1 _23066_ (.A1(_11173_),
    .A2(_11088_),
    .A3(_11185_),
    .A4(_11193_),
    .ZN(_13373_));
 NOR4_X1 _23067_ (.A1(_13371_),
    .A2(_13372_),
    .A3(_12647_),
    .A4(_13373_),
    .ZN(_13374_));
 AND4_X1 _23068_ (.A1(_13365_),
    .A2(_13367_),
    .A3(_13370_),
    .A4(_13374_),
    .ZN(_13375_));
 OAI21_X1 _23069_ (.A(_11234_),
    .B1(_12230_),
    .B2(_11225_),
    .ZN(_13376_));
 NAND2_X1 _23070_ (.A1(_12580_),
    .A2(_11252_),
    .ZN(_13377_));
 NAND2_X1 _23071_ (.A1(_11234_),
    .A2(_11105_),
    .ZN(_13378_));
 OAI21_X1 _23072_ (.A(_11252_),
    .B1(_11282_),
    .B2(_11248_),
    .ZN(_13379_));
 NAND4_X1 _23073_ (.A1(_13376_),
    .A2(_13377_),
    .A3(_13378_),
    .A4(_13379_),
    .ZN(_13380_));
 NAND4_X1 _23074_ (.A1(_11255_),
    .A2(_11238_),
    .A3(_11194_),
    .A4(_11155_),
    .ZN(_13381_));
 OAI221_X1 _23075_ (.A(_13381_),
    .B1(_12588_),
    .B2(_11111_),
    .C1(_11142_),
    .C2(_12279_),
    .ZN(_13382_));
 AOI21_X1 _23076_ (.A(_12588_),
    .B1(_12219_),
    .B2(_11218_),
    .ZN(_13383_));
 OAI21_X1 _23077_ (.A(_11247_),
    .B1(_12642_),
    .B2(_11304_),
    .ZN(_13384_));
 OAI21_X1 _23078_ (.A(_11247_),
    .B1(_11121_),
    .B2(_11139_),
    .ZN(_13385_));
 NAND2_X1 _23079_ (.A1(_11247_),
    .A2(_12226_),
    .ZN(_13386_));
 NAND4_X1 _23080_ (.A1(_13384_),
    .A2(_13385_),
    .A3(_11249_),
    .A4(_13386_),
    .ZN(_13387_));
 NOR4_X1 _23081_ (.A1(_13380_),
    .A2(_13382_),
    .A3(_13383_),
    .A4(_13387_),
    .ZN(_13388_));
 OAI21_X1 _23082_ (.A(_11285_),
    .B1(_11116_),
    .B2(_11121_),
    .ZN(_13389_));
 NAND2_X1 _23083_ (.A1(_11274_),
    .A2(_11110_),
    .ZN(_13390_));
 NAND4_X1 _23084_ (.A1(_11255_),
    .A2(_11194_),
    .A3(_11189_),
    .A4(_11288_),
    .ZN(_13391_));
 AND3_X1 _23085_ (.A1(_13389_),
    .A2(_13390_),
    .A3(_13391_),
    .ZN(_13392_));
 NAND2_X1 _23086_ (.A1(_11299_),
    .A2(_12830_),
    .ZN(_13393_));
 OAI21_X1 _23087_ (.A(_13393_),
    .B1(_12208_),
    .B2(_12202_),
    .ZN(_13394_));
 AND2_X1 _23088_ (.A1(_12275_),
    .A2(_11299_),
    .ZN(_13395_));
 AND3_X1 _23089_ (.A1(_11297_),
    .A2(_11115_),
    .A3(_11099_),
    .ZN(_13396_));
 NOR4_X1 _23090_ (.A1(_13394_),
    .A2(_13395_),
    .A3(_12207_),
    .A4(_13396_),
    .ZN(_13397_));
 AOI21_X1 _23091_ (.A(_12862_),
    .B1(_12251_),
    .B2(_11117_),
    .ZN(_13398_));
 AND2_X1 _23092_ (.A1(_12205_),
    .A2(_11264_),
    .ZN(_13399_));
 AND3_X1 _23093_ (.A1(_11181_),
    .A2(_12182_),
    .A3(_11288_),
    .ZN(_13400_));
 NOR4_X1 _23094_ (.A1(_13398_),
    .A2(_13176_),
    .A3(_13399_),
    .A4(_13400_),
    .ZN(_13401_));
 OAI21_X1 _23095_ (.A(_11295_),
    .B1(_11128_),
    .B2(_12822_),
    .ZN(_13402_));
 OAI21_X1 _23096_ (.A(_11295_),
    .B1(_11181_),
    .B2(_11160_),
    .ZN(_13403_));
 NAND4_X1 _23097_ (.A1(_11295_),
    .A2(_11184_),
    .A3(_11186_),
    .A4(_11194_),
    .ZN(_13404_));
 AND3_X1 _23098_ (.A1(_13402_),
    .A2(_13403_),
    .A3(_13404_),
    .ZN(_13405_));
 AND4_X1 _23099_ (.A1(_13392_),
    .A2(_13397_),
    .A3(_13401_),
    .A4(_13405_),
    .ZN(_13406_));
 NAND4_X1 _23100_ (.A1(_13361_),
    .A2(_13375_),
    .A3(_13388_),
    .A4(_13406_),
    .ZN(_13407_));
 NOR2_X2 _23101_ (.A1(_13407_),
    .A2(_11311_),
    .ZN(_13408_));
 AND4_X1 _23102_ (.A1(_11632_),
    .A2(_11616_),
    .A3(_11672_),
    .A4(_11637_),
    .ZN(_13409_));
 AOI221_X4 _23103_ (.A(_13409_),
    .B1(_11821_),
    .B2(_11577_),
    .C1(_12163_),
    .C2(_11824_),
    .ZN(_13410_));
 INV_X1 _23104_ (.A(_11782_),
    .ZN(_13411_));
 NAND3_X1 _23105_ (.A1(_11612_),
    .A2(_11572_),
    .A3(_11646_),
    .ZN(_13412_));
 OAI21_X1 _23106_ (.A(_11656_),
    .B1(_12112_),
    .B2(_11725_),
    .ZN(_13413_));
 OAI21_X1 _23107_ (.A(_11639_),
    .B1(_11622_),
    .B2(_11757_),
    .ZN(_13414_));
 AND4_X1 _23108_ (.A1(_13411_),
    .A2(_13412_),
    .A3(_13413_),
    .A4(_13414_),
    .ZN(_13415_));
 OAI21_X1 _23109_ (.A(_11821_),
    .B1(_11768_),
    .B2(_11644_),
    .ZN(_13416_));
 AOI21_X1 _23110_ (.A(_11818_),
    .B1(_11860_),
    .B2(_11746_),
    .ZN(_13417_));
 NAND2_X1 _23111_ (.A1(_11689_),
    .A2(_11667_),
    .ZN(_13418_));
 OAI21_X1 _23112_ (.A(_13418_),
    .B1(_11741_),
    .B2(_11818_),
    .ZN(_13419_));
 AND2_X1 _23113_ (.A1(_11833_),
    .A2(_11675_),
    .ZN(_13420_));
 NOR4_X1 _23114_ (.A1(_13417_),
    .A2(_13419_),
    .A3(_13420_),
    .A4(_11670_),
    .ZN(_13421_));
 AND4_X1 _23115_ (.A1(_13410_),
    .A2(_13415_),
    .A3(_13416_),
    .A4(_13421_),
    .ZN(_13422_));
 AOI221_X1 _23116_ (.A(_11717_),
    .B1(_11559_),
    .B2(_11582_),
    .C1(_11631_),
    .C2(_11786_),
    .ZN(_13423_));
 INV_X1 _23117_ (.A(_13138_),
    .ZN(_13424_));
 NOR4_X1 _23118_ (.A1(_13423_),
    .A2(_13424_),
    .A3(_12130_),
    .A4(_12131_),
    .ZN(_13425_));
 OAI21_X1 _23119_ (.A(_11680_),
    .B1(_12171_),
    .B2(_11761_),
    .ZN(_13426_));
 AND3_X1 _23120_ (.A1(_13426_),
    .A2(_11855_),
    .A3(_13136_),
    .ZN(_13427_));
 NAND2_X1 _23121_ (.A1(_11722_),
    .A2(_11799_),
    .ZN(_13428_));
 OAI21_X1 _23122_ (.A(_11722_),
    .B1(_11720_),
    .B2(_12529_),
    .ZN(_13429_));
 NAND2_X1 _23123_ (.A1(_11722_),
    .A2(_11768_),
    .ZN(_13430_));
 AND4_X1 _23124_ (.A1(_13428_),
    .A2(_13429_),
    .A3(_13430_),
    .A4(_12537_),
    .ZN(_13431_));
 AND2_X1 _23125_ (.A1(_11587_),
    .A2(_11704_),
    .ZN(_13432_));
 AOI211_X1 _23126_ (.A(_11697_),
    .B(_13432_),
    .C1(_11705_),
    .C2(_11704_),
    .ZN(_13433_));
 AND4_X1 _23127_ (.A1(_13425_),
    .A2(_13427_),
    .A3(_13431_),
    .A4(_13433_),
    .ZN(_13434_));
 OAI21_X1 _23128_ (.A(_11607_),
    .B1(_11683_),
    .B2(_11622_),
    .ZN(_13435_));
 OAI21_X1 _23129_ (.A(_11607_),
    .B1(_11689_),
    .B2(_11768_),
    .ZN(_13436_));
 AND3_X1 _23130_ (.A1(_13435_),
    .A2(_13436_),
    .A3(_11613_),
    .ZN(_13437_));
 NAND3_X1 _23131_ (.A1(_11627_),
    .A2(_11588_),
    .A3(_11566_),
    .ZN(_13438_));
 OAI21_X1 _23132_ (.A(_11581_),
    .B1(_11737_),
    .B2(_11587_),
    .ZN(_13439_));
 AND4_X1 _23133_ (.A1(_11585_),
    .A2(_13127_),
    .A3(_13438_),
    .A4(_13439_),
    .ZN(_13440_));
 INV_X1 _23134_ (.A(_12510_),
    .ZN(_13441_));
 NAND3_X1 _23135_ (.A1(_12149_),
    .A2(_11706_),
    .A3(_16698_),
    .ZN(_13442_));
 AND4_X1 _23136_ (.A1(_13441_),
    .A2(_11837_),
    .A3(_13132_),
    .A4(_13442_),
    .ZN(_13443_));
 OAI21_X1 _23137_ (.A(_11553_),
    .B1(_11694_),
    .B2(_11598_),
    .ZN(_13444_));
 AND3_X1 _23138_ (.A1(_13444_),
    .A2(_11565_),
    .A3(_11573_),
    .ZN(_13445_));
 AND4_X1 _23139_ (.A1(_13437_),
    .A2(_13440_),
    .A3(_13443_),
    .A4(_13445_),
    .ZN(_13446_));
 OAI21_X1 _23140_ (.A(_12122_),
    .B1(_12506_),
    .B2(_12938_),
    .ZN(_13447_));
 OAI21_X1 _23141_ (.A(_12122_),
    .B1(_11687_),
    .B2(_11577_),
    .ZN(_13448_));
 OAI211_X1 _23142_ (.A(_12122_),
    .B(_11702_),
    .C1(_11701_),
    .C2(_11661_),
    .ZN(_13449_));
 AND3_X1 _23143_ (.A1(_13447_),
    .A2(_13448_),
    .A3(_13449_),
    .ZN(_13450_));
 OAI211_X1 _23144_ (.A(_11735_),
    .B(_11709_),
    .C1(_11706_),
    .C2(_11707_),
    .ZN(_13451_));
 AND4_X1 _23145_ (.A1(_13121_),
    .A2(_13122_),
    .A3(_12571_),
    .A4(_13451_),
    .ZN(_13452_));
 NOR2_X1 _23146_ (.A1(_12504_),
    .A2(_12116_),
    .ZN(_13453_));
 AND2_X1 _23147_ (.A1(_11756_),
    .A2(_11577_),
    .ZN(_13454_));
 AND4_X1 _23148_ (.A1(_11732_),
    .A2(_11659_),
    .A3(_11672_),
    .A4(_11710_),
    .ZN(_13455_));
 NOR3_X1 _23149_ (.A1(_13453_),
    .A2(_13454_),
    .A3(_13455_),
    .ZN(_13456_));
 NAND3_X1 _23150_ (.A1(_11767_),
    .A2(_11661_),
    .A3(_11592_),
    .ZN(_13457_));
 OAI211_X1 _23151_ (.A(_11767_),
    .B(_11702_),
    .C1(_11706_),
    .C2(_11707_),
    .ZN(_13458_));
 NAND4_X1 _23152_ (.A1(_11709_),
    .A2(_11701_),
    .A3(_11732_),
    .A4(_11588_),
    .ZN(_13459_));
 AND4_X1 _23153_ (.A1(_13457_),
    .A2(_13458_),
    .A3(_11800_),
    .A4(_13459_),
    .ZN(_13460_));
 AND4_X1 _23154_ (.A1(_13450_),
    .A2(_13452_),
    .A3(_13456_),
    .A4(_13460_),
    .ZN(_13461_));
 NAND4_X1 _23155_ (.A1(_13422_),
    .A2(_13434_),
    .A3(_13446_),
    .A4(_13461_),
    .ZN(_13462_));
 NOR2_X2 _23156_ (.A1(_13462_),
    .A2(_11775_),
    .ZN(_13463_));
 XNOR2_X2 _23157_ (.A(_13408_),
    .B(_13463_),
    .ZN(_13464_));
 OAI21_X1 _23158_ (.A(_12094_),
    .B1(_11964_),
    .B2(_12027_),
    .ZN(_13465_));
 AND2_X1 _23159_ (.A1(_11948_),
    .A2(_12088_),
    .ZN(_13466_));
 AND2_X1 _23160_ (.A1(_11929_),
    .A2(_12089_),
    .ZN(_13467_));
 AOI211_X1 _23161_ (.A(_13466_),
    .B(_13467_),
    .C1(_12089_),
    .C2(_12014_),
    .ZN(_13468_));
 OAI211_X1 _23162_ (.A(_12094_),
    .B(_12397_),
    .C1(_11955_),
    .C2(_12414_),
    .ZN(_13469_));
 OAI21_X1 _23163_ (.A(_12094_),
    .B1(_12024_),
    .B2(_12412_),
    .ZN(_13470_));
 AND4_X1 _23164_ (.A1(_13465_),
    .A2(_13468_),
    .A3(_13469_),
    .A4(_13470_),
    .ZN(_13471_));
 NAND2_X1 _23165_ (.A1(_11989_),
    .A2(_12423_),
    .ZN(_13472_));
 NAND2_X1 _23166_ (.A1(_12737_),
    .A2(_12064_),
    .ZN(_13473_));
 OAI211_X1 _23167_ (.A(_12423_),
    .B(_12011_),
    .C1(_11932_),
    .C2(_11933_),
    .ZN(_13474_));
 NAND4_X1 _23168_ (.A1(_13472_),
    .A2(_13273_),
    .A3(_13473_),
    .A4(_13474_),
    .ZN(_13475_));
 AOI211_X1 _23169_ (.A(_11916_),
    .B(_12445_),
    .C1(_11880_),
    .C2(_11919_),
    .ZN(_13476_));
 NAND2_X1 _23170_ (.A1(_12440_),
    .A2(_12455_),
    .ZN(_13477_));
 OAI22_X1 _23171_ (.A1(_13477_),
    .A2(_11946_),
    .B1(_12445_),
    .B2(_12013_),
    .ZN(_13478_));
 NOR3_X1 _23172_ (.A1(_13475_),
    .A2(_13476_),
    .A3(_13478_),
    .ZN(_13479_));
 OAI211_X1 _23173_ (.A(_12073_),
    .B(_12428_),
    .C1(_12069_),
    .C2(_12432_),
    .ZN(_13480_));
 AOI21_X1 _23174_ (.A(_12069_),
    .B1(_12083_),
    .B2(_12743_),
    .ZN(_13481_));
 AOI21_X1 _23175_ (.A(_12079_),
    .B1(_11986_),
    .B2(_12781_),
    .ZN(_13482_));
 NOR4_X1 _23176_ (.A1(_13480_),
    .A2(_13481_),
    .A3(_13482_),
    .A4(_12788_),
    .ZN(_13483_));
 AND2_X1 _23177_ (.A1(_12027_),
    .A2(_12030_),
    .ZN(_13484_));
 INV_X1 _23178_ (.A(_13484_),
    .ZN(_13485_));
 NAND2_X1 _23179_ (.A1(_12022_),
    .A2(_11929_),
    .ZN(_13486_));
 OAI21_X1 _23180_ (.A(_12022_),
    .B1(_12033_),
    .B2(_11937_),
    .ZN(_13487_));
 OAI21_X1 _23181_ (.A(_12022_),
    .B1(_12003_),
    .B2(_12410_),
    .ZN(_13488_));
 NAND2_X1 _23182_ (.A1(_12019_),
    .A2(_12447_),
    .ZN(_13489_));
 AND4_X1 _23183_ (.A1(_13486_),
    .A2(_13487_),
    .A3(_13488_),
    .A4(_13489_),
    .ZN(_13490_));
 OAI21_X1 _23184_ (.A(_12391_),
    .B1(_12417_),
    .B2(_12034_),
    .ZN(_13491_));
 AND4_X1 _23185_ (.A1(_13485_),
    .A2(_13490_),
    .A3(_13010_),
    .A4(_13491_),
    .ZN(_13492_));
 NAND4_X1 _23186_ (.A1(_13471_),
    .A2(_13479_),
    .A3(_13483_),
    .A4(_13492_),
    .ZN(_13493_));
 AOI22_X1 _23187_ (.A1(_12801_),
    .A2(_12429_),
    .B1(_12090_),
    .B2(_11974_),
    .ZN(_13494_));
 OAI21_X1 _23188_ (.A(_11993_),
    .B1(_12055_),
    .B2(_12090_),
    .ZN(_13495_));
 OAI21_X1 _23189_ (.A(_11974_),
    .B1(_12737_),
    .B2(_12447_),
    .ZN(_13496_));
 AND4_X1 _23190_ (.A1(_12771_),
    .A2(_13494_),
    .A3(_13495_),
    .A4(_13496_),
    .ZN(_13497_));
 NAND2_X1 _23191_ (.A1(_12480_),
    .A2(_11900_),
    .ZN(_13498_));
 NAND3_X1 _23192_ (.A1(_11960_),
    .A2(_11963_),
    .A3(_13498_),
    .ZN(_13499_));
 NAND2_X1 _23193_ (.A1(_12480_),
    .A2(_11929_),
    .ZN(_13500_));
 OAI211_X1 _23194_ (.A(_13500_),
    .B(_13219_),
    .C1(_12481_),
    .C2(_12083_),
    .ZN(_13501_));
 AOI21_X1 _23195_ (.A(_12753_),
    .B1(_12781_),
    .B2(_12432_),
    .ZN(_13502_));
 NOR4_X1 _23196_ (.A1(_13499_),
    .A2(_13501_),
    .A3(_12973_),
    .A4(_13502_),
    .ZN(_13503_));
 OAI21_X1 _23197_ (.A(_12762_),
    .B1(_12417_),
    .B2(_12449_),
    .ZN(_13504_));
 OAI211_X1 _23198_ (.A(_12489_),
    .B(_16786_),
    .C1(_16785_),
    .C2(_11927_),
    .ZN(_13505_));
 OAI21_X1 _23199_ (.A(_12762_),
    .B1(_11994_),
    .B2(_12084_),
    .ZN(_13506_));
 AND4_X1 _23200_ (.A1(_12488_),
    .A2(_13504_),
    .A3(_13505_),
    .A4(_13506_),
    .ZN(_13507_));
 AND2_X1 _23201_ (.A1(_12465_),
    .A2(_12466_),
    .ZN(_13508_));
 NAND3_X1 _23202_ (.A1(_11894_),
    .A2(_11911_),
    .A3(_11979_),
    .ZN(_13509_));
 AND3_X1 _23203_ (.A1(_12739_),
    .A2(_13236_),
    .A3(_13509_),
    .ZN(_13510_));
 OAI21_X1 _23204_ (.A(_12461_),
    .B1(_11898_),
    .B2(_11894_),
    .ZN(_13511_));
 OAI21_X1 _23205_ (.A(_12461_),
    .B1(_11970_),
    .B2(_11953_),
    .ZN(_13512_));
 AND4_X1 _23206_ (.A1(_13508_),
    .A2(_13510_),
    .A3(_13511_),
    .A4(_13512_),
    .ZN(_13513_));
 NAND4_X1 _23207_ (.A1(_13497_),
    .A2(_13503_),
    .A3(_13507_),
    .A4(_13513_),
    .ZN(_13514_));
 NOR2_X2 _23208_ (.A1(_13493_),
    .A2(_13514_),
    .ZN(_13515_));
 XOR2_X2 _23209_ (.A(_13464_),
    .B(_13515_),
    .Z(_13516_));
 AND2_X1 _23210_ (.A1(_11425_),
    .A2(_11487_),
    .ZN(_13517_));
 OR3_X1 _23211_ (.A1(_13045_),
    .A2(_12667_),
    .A3(_13517_),
    .ZN(_13518_));
 OR3_X1 _23212_ (.A1(_11471_),
    .A2(_11514_),
    .A3(_11509_),
    .ZN(_13519_));
 AOI22_X1 _23213_ (.A1(_11410_),
    .A2(_12366_),
    .B1(_11536_),
    .B2(_12322_),
    .ZN(_13520_));
 OAI211_X1 _23214_ (.A(_13520_),
    .B(_12662_),
    .C1(_11526_),
    .C2(_11387_),
    .ZN(_13521_));
 OAI211_X1 _23215_ (.A(_12678_),
    .B(_12294_),
    .C1(_12345_),
    .C2(_11390_),
    .ZN(_13522_));
 NOR4_X1 _23216_ (.A1(_13518_),
    .A2(_13519_),
    .A3(_13521_),
    .A4(_13522_),
    .ZN(_13523_));
 AOI21_X1 _23217_ (.A(_12697_),
    .B1(_11341_),
    .B2(_12346_),
    .ZN(_13524_));
 AND2_X1 _23218_ (.A1(_12375_),
    .A2(_11406_),
    .ZN(_13525_));
 NOR3_X1 _23219_ (.A1(_13524_),
    .A2(_11455_),
    .A3(_13525_),
    .ZN(_13526_));
 AND2_X1 _23220_ (.A1(_11477_),
    .A2(_11442_),
    .ZN(_13527_));
 AND3_X1 _23221_ (.A1(_12321_),
    .A2(_11381_),
    .A3(_11349_),
    .ZN(_13528_));
 AND3_X1 _23222_ (.A1(_11442_),
    .A2(_11316_),
    .A3(_11349_),
    .ZN(_13529_));
 NOR4_X1 _23223_ (.A1(_12652_),
    .A2(_13527_),
    .A3(_13528_),
    .A4(_13529_),
    .ZN(_13530_));
 NAND2_X1 _23224_ (.A1(_11434_),
    .A2(_11398_),
    .ZN(_13531_));
 OAI21_X1 _23225_ (.A(_11414_),
    .B1(_11511_),
    .B2(_11461_),
    .ZN(_13532_));
 NAND3_X1 _23226_ (.A1(_12337_),
    .A2(_11534_),
    .A3(_11472_),
    .ZN(_13533_));
 NAND2_X1 _23227_ (.A1(_11493_),
    .A2(_11405_),
    .ZN(_13534_));
 AND4_X1 _23228_ (.A1(_13531_),
    .A2(_13532_),
    .A3(_13533_),
    .A4(_13534_),
    .ZN(_13535_));
 NAND2_X1 _23229_ (.A1(_11420_),
    .A2(_11450_),
    .ZN(_13536_));
 OAI21_X1 _23230_ (.A(_13536_),
    .B1(_13305_),
    .B2(_12288_),
    .ZN(_13537_));
 AND3_X1 _23231_ (.A1(_11356_),
    .A2(_11534_),
    .A3(_11408_),
    .ZN(_13538_));
 NOR2_X1 _23232_ (.A1(_13537_),
    .A2(_13538_),
    .ZN(_13539_));
 AND4_X1 _23233_ (.A1(_13526_),
    .A2(_13530_),
    .A3(_13535_),
    .A4(_13539_),
    .ZN(_13540_));
 NAND2_X1 _23234_ (.A1(_11518_),
    .A2(_11406_),
    .ZN(_13541_));
 OAI21_X1 _23235_ (.A(_11488_),
    .B1(_11363_),
    .B2(_11542_),
    .ZN(_13542_));
 OAI21_X1 _23236_ (.A(_11482_),
    .B1(_11373_),
    .B2(_13084_),
    .ZN(_13543_));
 OAI21_X1 _23237_ (.A(_11434_),
    .B1(_11410_),
    .B2(_11452_),
    .ZN(_13544_));
 AND4_X1 _23238_ (.A1(_13541_),
    .A2(_13542_),
    .A3(_13543_),
    .A4(_13544_),
    .ZN(_13545_));
 NAND2_X1 _23239_ (.A1(_12366_),
    .A2(_11511_),
    .ZN(_13546_));
 NAND3_X1 _23240_ (.A1(_12371_),
    .A2(_13546_),
    .A3(_13328_),
    .ZN(_13547_));
 NOR2_X1 _23241_ (.A1(_13315_),
    .A2(_11362_),
    .ZN(_13548_));
 AND2_X1 _23242_ (.A1(_11467_),
    .A2(_11459_),
    .ZN(_13549_));
 AND2_X1 _23243_ (.A1(_11366_),
    .A2(_11326_),
    .ZN(_13550_));
 NOR4_X1 _23244_ (.A1(_13547_),
    .A2(_13548_),
    .A3(_13549_),
    .A4(_13550_),
    .ZN(_13551_));
 NAND4_X1 _23245_ (.A1(_13523_),
    .A2(_13540_),
    .A3(_13545_),
    .A4(_13551_),
    .ZN(_13552_));
 AND2_X1 _23246_ (.A1(_11522_),
    .A2(_11437_),
    .ZN(_13553_));
 AND2_X1 _23247_ (.A1(_11542_),
    .A2(_11481_),
    .ZN(_13554_));
 AND2_X1 _23248_ (.A1(_11382_),
    .A2(_11344_),
    .ZN(_13555_));
 AND2_X1 _23249_ (.A1(_11410_),
    .A2(_11386_),
    .ZN(_13556_));
 NOR4_X1 _23250_ (.A1(_13553_),
    .A2(_13554_),
    .A3(_13555_),
    .A4(_13556_),
    .ZN(_13557_));
 INV_X1 _23251_ (.A(_13031_),
    .ZN(_13558_));
 AOI22_X1 _23252_ (.A1(_11482_),
    .A2(_12690_),
    .B1(_12375_),
    .B2(_11431_),
    .ZN(_13559_));
 AND4_X1 _23253_ (.A1(_11337_),
    .A2(_13557_),
    .A3(_13558_),
    .A4(_13559_),
    .ZN(_13560_));
 AND2_X1 _23254_ (.A1(_11511_),
    .A2(_11318_),
    .ZN(_13561_));
 AOI211_X1 _23255_ (.A(_11322_),
    .B(_13561_),
    .C1(_11403_),
    .C2(_11437_),
    .ZN(_13562_));
 OAI211_X1 _23256_ (.A(_11403_),
    .B(_11373_),
    .C1(_11338_),
    .C2(_11472_),
    .ZN(_13563_));
 AND3_X1 _23257_ (.A1(_11352_),
    .A2(_13036_),
    .A3(_12664_),
    .ZN(_13564_));
 AND4_X1 _23258_ (.A1(_11362_),
    .A2(_11368_),
    .A3(_11351_),
    .A4(_11334_),
    .ZN(_13565_));
 NOR3_X1 _23259_ (.A1(_13564_),
    .A2(_12669_),
    .A3(_13565_),
    .ZN(_13566_));
 OAI21_X1 _23260_ (.A(_11431_),
    .B1(_11540_),
    .B2(_13070_),
    .ZN(_13567_));
 AND4_X1 _23261_ (.A1(_13562_),
    .A2(_13563_),
    .A3(_13566_),
    .A4(_13567_),
    .ZN(_13568_));
 INV_X1 _23262_ (.A(_11449_),
    .ZN(_13569_));
 AND4_X1 _23263_ (.A1(_13312_),
    .A2(_11500_),
    .A3(_13057_),
    .A4(_13313_),
    .ZN(_13570_));
 NAND2_X1 _23264_ (.A1(_11347_),
    .A2(_11456_),
    .ZN(_13571_));
 OAI21_X1 _23265_ (.A(_11525_),
    .B1(_12366_),
    .B2(_11488_),
    .ZN(_13572_));
 AND4_X1 _23266_ (.A1(_13569_),
    .A2(_13570_),
    .A3(_13571_),
    .A4(_13572_),
    .ZN(_13573_));
 AOI22_X1 _23267_ (.A1(_12338_),
    .A2(_11415_),
    .B1(_11460_),
    .B2(_13084_),
    .ZN(_13574_));
 AOI22_X1 _23268_ (.A1(_11467_),
    .A2(_12374_),
    .B1(_11410_),
    .B2(_11415_),
    .ZN(_13575_));
 AOI22_X1 _23269_ (.A1(_11353_),
    .A2(_11321_),
    .B1(_11420_),
    .B2(_11483_),
    .ZN(_13576_));
 AOI22_X1 _23270_ (.A1(_12296_),
    .A2(_11460_),
    .B1(_11414_),
    .B2(_11327_),
    .ZN(_13577_));
 AND4_X1 _23271_ (.A1(_13574_),
    .A2(_13575_),
    .A3(_13576_),
    .A4(_13577_),
    .ZN(_13578_));
 NAND4_X1 _23272_ (.A1(_13560_),
    .A2(_13568_),
    .A3(_13573_),
    .A4(_13578_),
    .ZN(_13579_));
 NOR2_X2 _23273_ (.A1(_13552_),
    .A2(_13579_),
    .ZN(_13580_));
 XOR2_X1 _23274_ (.A(_13159_),
    .B(_13580_),
    .Z(_13581_));
 XNOR2_X1 _23275_ (.A(_13516_),
    .B(_13581_),
    .ZN(_13582_));
 XNOR2_X1 _23276_ (.A(_13582_),
    .B(_17190_),
    .ZN(_13583_));
 MUX2_X1 _23277_ (.A(_13350_),
    .B(_13583_),
    .S(_11084_),
    .Z(_00721_));
 XOR2_X1 _23278_ (.A(_17191_),
    .B(_16994_),
    .Z(_13584_));
 OAI21_X1 _23279_ (.A(_11265_),
    .B1(_11128_),
    .B2(_12822_),
    .ZN(_13585_));
 NAND3_X1 _23280_ (.A1(_11265_),
    .A2(_12239_),
    .A3(_11270_),
    .ZN(_13586_));
 NAND4_X1 _23281_ (.A1(_11194_),
    .A2(_12182_),
    .A3(_11173_),
    .A4(_11288_),
    .ZN(_13587_));
 AND3_X1 _23282_ (.A1(_13585_),
    .A2(_13586_),
    .A3(_13587_),
    .ZN(_13588_));
 NAND4_X1 _23283_ (.A1(_11137_),
    .A2(_11184_),
    .A3(_11186_),
    .A4(_11100_),
    .ZN(_13589_));
 OAI21_X1 _23284_ (.A(_11137_),
    .B1(_11128_),
    .B2(_12822_),
    .ZN(_13590_));
 AND3_X1 _23285_ (.A1(_13588_),
    .A2(_13589_),
    .A3(_13590_),
    .ZN(_13591_));
 OAI22_X1 _23286_ (.A1(_12218_),
    .A2(_12623_),
    .B1(_11117_),
    .B2(_12250_),
    .ZN(_13592_));
 NOR4_X1 _23287_ (.A1(_13592_),
    .A2(_12271_),
    .A3(_11198_),
    .A4(_12195_),
    .ZN(_13593_));
 OAI22_X1 _23288_ (.A1(_12588_),
    .A2(_11278_),
    .B1(_11107_),
    .B2(_12202_),
    .ZN(_13594_));
 AOI211_X1 _23289_ (.A(_12234_),
    .B(_13594_),
    .C1(_11166_),
    .C2(_11093_),
    .ZN(_13595_));
 AOI22_X1 _23290_ (.A1(_11252_),
    .A2(_11248_),
    .B1(_11149_),
    .B2(_11156_),
    .ZN(_13596_));
 NAND3_X1 _23291_ (.A1(_11116_),
    .A2(_11255_),
    .A3(_11288_),
    .ZN(_13597_));
 AOI22_X1 _23292_ (.A1(_11302_),
    .A2(_11251_),
    .B1(_11213_),
    .B2(_11304_),
    .ZN(_13598_));
 AOI22_X1 _23293_ (.A1(_11213_),
    .A2(_12275_),
    .B1(_11215_),
    .B2(_11191_),
    .ZN(_13599_));
 AOI22_X1 _23294_ (.A1(_11282_),
    .A2(_11274_),
    .B1(_11148_),
    .B2(_11301_),
    .ZN(_13600_));
 AND4_X1 _23295_ (.A1(_13597_),
    .A2(_13598_),
    .A3(_13599_),
    .A4(_13600_),
    .ZN(_13601_));
 AND4_X1 _23296_ (.A1(_13593_),
    .A2(_13595_),
    .A3(_13596_),
    .A4(_13601_),
    .ZN(_13602_));
 INV_X1 _23297_ (.A(_11311_),
    .ZN(_13603_));
 OAI211_X1 _23298_ (.A(_11247_),
    .B(_16738_),
    .C1(_11109_),
    .C2(_11097_),
    .ZN(_13604_));
 OAI211_X1 _23299_ (.A(_11237_),
    .B(_11195_),
    .C1(_11105_),
    .C2(_11160_),
    .ZN(_13605_));
 OAI21_X1 _23300_ (.A(_11247_),
    .B1(_12205_),
    .B2(_11177_),
    .ZN(_13606_));
 AND4_X1 _23301_ (.A1(_13603_),
    .A2(_13604_),
    .A3(_13605_),
    .A4(_13606_),
    .ZN(_13607_));
 OAI21_X1 _23302_ (.A(_11207_),
    .B1(_11152_),
    .B2(_11282_),
    .ZN(_13608_));
 OAI21_X1 _23303_ (.A(_11207_),
    .B1(_12829_),
    .B2(_11235_),
    .ZN(_13609_));
 AND4_X1 _23304_ (.A1(_12815_),
    .A2(_13607_),
    .A3(_13608_),
    .A4(_13609_),
    .ZN(_13610_));
 AND2_X1 _23305_ (.A1(_12605_),
    .A2(_12836_),
    .ZN(_13611_));
 AOI22_X1 _23306_ (.A1(_12864_),
    .A2(_11259_),
    .B1(_11139_),
    .B2(_11221_),
    .ZN(_13612_));
 AOI22_X1 _23307_ (.A1(_11279_),
    .A2(_11093_),
    .B1(_11302_),
    .B2(_11295_),
    .ZN(_13613_));
 AOI22_X1 _23308_ (.A1(_11152_),
    .A2(_11221_),
    .B1(_11234_),
    .B2(_11139_),
    .ZN(_13614_));
 AND4_X1 _23309_ (.A1(_13611_),
    .A2(_13612_),
    .A3(_13613_),
    .A4(_13614_),
    .ZN(_13615_));
 AND4_X1 _23310_ (.A1(_13591_),
    .A2(_13602_),
    .A3(_13610_),
    .A4(_13615_),
    .ZN(_13616_));
 NAND2_X1 _23311_ (.A1(_12623_),
    .A2(_12227_),
    .ZN(_13617_));
 OAI21_X1 _23312_ (.A(_11295_),
    .B1(_13617_),
    .B2(_12187_),
    .ZN(_13618_));
 NAND4_X1 _23313_ (.A1(_11091_),
    .A2(_11173_),
    .A3(_11195_),
    .A4(_11239_),
    .ZN(_13619_));
 NAND2_X1 _23314_ (.A1(_12226_),
    .A2(_11129_),
    .ZN(_13620_));
 OAI21_X1 _23315_ (.A(_11092_),
    .B1(_11282_),
    .B2(_11215_),
    .ZN(_13621_));
 NAND4_X1 _23316_ (.A1(_13618_),
    .A2(_13619_),
    .A3(_13620_),
    .A4(_13621_),
    .ZN(_13622_));
 AND2_X1 _23317_ (.A1(_11285_),
    .A2(_12199_),
    .ZN(_13623_));
 OR4_X1 _23318_ (.A1(_12277_),
    .A2(_13622_),
    .A3(_13623_),
    .A4(_13160_),
    .ZN(_13624_));
 OAI21_X1 _23319_ (.A(_11234_),
    .B1(_12221_),
    .B2(_12822_),
    .ZN(_13625_));
 OAI21_X1 _23320_ (.A(_13625_),
    .B1(_12198_),
    .B2(_12224_),
    .ZN(_13626_));
 OAI21_X1 _23321_ (.A(_11299_),
    .B1(_12642_),
    .B2(_11128_),
    .ZN(_13627_));
 OAI211_X1 _23322_ (.A(_11299_),
    .B(_11100_),
    .C1(_11150_),
    .C2(_11142_),
    .ZN(_13628_));
 OAI211_X1 _23323_ (.A(_13627_),
    .B(_13628_),
    .C1(_11172_),
    .C2(_12631_),
    .ZN(_13629_));
 AND3_X1 _23324_ (.A1(_11234_),
    .A2(_12239_),
    .A3(_11270_),
    .ZN(_13630_));
 AND2_X1 _23325_ (.A1(_11199_),
    .A2(_11096_),
    .ZN(_13631_));
 NOR2_X1 _23326_ (.A1(_13630_),
    .A2(_13631_),
    .ZN(_13632_));
 NAND3_X1 _23327_ (.A1(_11100_),
    .A2(_11193_),
    .A3(_11143_),
    .ZN(_13633_));
 AOI22_X1 _23328_ (.A1(_11259_),
    .A2(_11235_),
    .B1(_11285_),
    .B2(_11160_),
    .ZN(_13634_));
 NAND4_X1 _23329_ (.A1(_13632_),
    .A2(_12632_),
    .A3(_13633_),
    .A4(_13634_),
    .ZN(_13635_));
 NOR4_X1 _23330_ (.A1(_13624_),
    .A2(_13626_),
    .A3(_13629_),
    .A4(_13635_),
    .ZN(_13636_));
 AND2_X1 _23331_ (.A1(_13616_),
    .A2(_13636_),
    .ZN(_13637_));
 NOR3_X1 _23332_ (.A1(_11665_),
    .A2(_11822_),
    .A3(_12888_),
    .ZN(_13638_));
 INV_X1 _23333_ (.A(_12164_),
    .ZN(_13639_));
 OAI211_X1 _23334_ (.A(_13638_),
    .B(_13639_),
    .C1(_12544_),
    .C2(_11840_),
    .ZN(_13640_));
 AND2_X1 _23335_ (.A1(_11759_),
    .A2(_11656_),
    .ZN(_13641_));
 OAI21_X1 _23336_ (.A(_12169_),
    .B1(_11652_),
    .B2(_11746_),
    .ZN(_13642_));
 AND4_X1 _23337_ (.A1(_11824_),
    .A2(_11672_),
    .A3(_11646_),
    .A4(_11572_),
    .ZN(_13643_));
 AND4_X1 _23338_ (.A1(_11824_),
    .A2(_11571_),
    .A3(_11646_),
    .A4(_11572_),
    .ZN(_13644_));
 OR4_X1 _23339_ (.A1(_13641_),
    .A2(_13642_),
    .A3(_13643_),
    .A4(_13644_),
    .ZN(_13645_));
 OAI211_X1 _23340_ (.A(_11675_),
    .B(_11702_),
    .C1(_11701_),
    .C2(_11661_),
    .ZN(_13646_));
 OAI211_X1 _23341_ (.A(_11675_),
    .B(_16698_),
    .C1(_11707_),
    .C2(_11554_),
    .ZN(_13647_));
 OAI21_X1 _23342_ (.A(_11675_),
    .B1(_11612_),
    .B2(_11577_),
    .ZN(_13648_));
 NAND3_X1 _23343_ (.A1(_13646_),
    .A2(_13647_),
    .A3(_13648_),
    .ZN(_13649_));
 OAI21_X1 _23344_ (.A(_11639_),
    .B1(_11687_),
    .B2(_11757_),
    .ZN(_13650_));
 OAI211_X1 _23345_ (.A(_13650_),
    .B(_12177_),
    .C1(_11783_),
    .C2(_11796_),
    .ZN(_13651_));
 NOR4_X1 _23346_ (.A1(_13640_),
    .A2(_13645_),
    .A3(_13649_),
    .A4(_13651_),
    .ZN(_13652_));
 AND2_X1 _23347_ (.A1(_12149_),
    .A2(_11622_),
    .ZN(_13653_));
 AOI21_X1 _23348_ (.A(_11618_),
    .B1(_11594_),
    .B2(_11595_),
    .ZN(_13654_));
 AND3_X1 _23349_ (.A1(_11674_),
    .A2(_11566_),
    .A3(_11616_),
    .ZN(_13655_));
 OR4_X1 _23350_ (.A1(_13653_),
    .A2(_13654_),
    .A3(_11634_),
    .A4(_13655_),
    .ZN(_13656_));
 OAI21_X1 _23351_ (.A(_11553_),
    .B1(_12506_),
    .B2(_12938_),
    .ZN(_13657_));
 OAI21_X1 _23352_ (.A(_13657_),
    .B1(_12533_),
    .B2(_11847_),
    .ZN(_13658_));
 OAI21_X1 _23353_ (.A(_11607_),
    .B1(_11598_),
    .B2(_12529_),
    .ZN(_13659_));
 OAI211_X1 _23354_ (.A(_13659_),
    .B(_12920_),
    .C1(_11811_),
    .C2(_11843_),
    .ZN(_13660_));
 OAI21_X1 _23355_ (.A(_11834_),
    .B1(_11591_),
    .B2(_11654_),
    .ZN(_13661_));
 OR3_X1 _23356_ (.A1(_13661_),
    .A2(_11830_),
    .A3(_11831_),
    .ZN(_13662_));
 NOR4_X1 _23357_ (.A1(_13656_),
    .A2(_13658_),
    .A3(_13660_),
    .A4(_13662_),
    .ZN(_13663_));
 NOR4_X1 _23358_ (.A1(_12525_),
    .A2(_12526_),
    .A3(_13424_),
    .A4(_12130_),
    .ZN(_13664_));
 NAND2_X1 _23359_ (.A1(_11722_),
    .A2(_11564_),
    .ZN(_13665_));
 AND4_X1 _23360_ (.A1(_13430_),
    .A2(_11866_),
    .A3(_13665_),
    .A4(_12946_),
    .ZN(_13666_));
 AOI21_X1 _23361_ (.A(_11692_),
    .B1(_11778_),
    .B2(_11840_),
    .ZN(_13667_));
 AND4_X1 _23362_ (.A1(_11642_),
    .A2(_11602_),
    .A3(_11672_),
    .A4(_11695_),
    .ZN(_13668_));
 NOR4_X1 _23363_ (.A1(_13667_),
    .A2(_12934_),
    .A3(_12935_),
    .A4(_13668_),
    .ZN(_13669_));
 AND2_X1 _23364_ (.A1(_11609_),
    .A2(_11704_),
    .ZN(_13670_));
 NOR4_X1 _23365_ (.A1(_13670_),
    .A2(_13432_),
    .A3(_12949_),
    .A4(_11699_),
    .ZN(_13671_));
 AND4_X1 _23366_ (.A1(_13664_),
    .A2(_13666_),
    .A3(_13669_),
    .A4(_13671_),
    .ZN(_13672_));
 OAI21_X1 _23367_ (.A(_11735_),
    .B1(_12506_),
    .B2(_12938_),
    .ZN(_13673_));
 NAND3_X1 _23368_ (.A1(_11735_),
    .A2(_11669_),
    .A3(_11671_),
    .ZN(_13674_));
 NAND4_X1 _23369_ (.A1(_11602_),
    .A2(_11702_),
    .A3(_11824_),
    .A4(_11732_),
    .ZN(_13675_));
 AND3_X1 _23370_ (.A1(_13673_),
    .A2(_13674_),
    .A3(_13675_),
    .ZN(_13676_));
 AOI21_X1 _23371_ (.A(_12116_),
    .B1(_11691_),
    .B2(_11796_),
    .ZN(_13677_));
 NOR3_X1 _23372_ (.A1(_13677_),
    .A2(_12897_),
    .A3(_13454_),
    .ZN(_13678_));
 AOI21_X1 _23373_ (.A(_11747_),
    .B1(_11628_),
    .B2(_11848_),
    .ZN(_13679_));
 AOI21_X1 _23374_ (.A(_11747_),
    .B1(_11780_),
    .B2(_11811_),
    .ZN(_13680_));
 NOR3_X1 _23375_ (.A1(_13679_),
    .A2(_13680_),
    .A3(_12124_),
    .ZN(_13681_));
 OAI21_X1 _23376_ (.A(_11767_),
    .B1(_12508_),
    .B2(_11809_),
    .ZN(_13682_));
 AND4_X1 _23377_ (.A1(_13676_),
    .A2(_13678_),
    .A3(_13681_),
    .A4(_13682_),
    .ZN(_13683_));
 NAND4_X1 _23378_ (.A1(_13652_),
    .A2(_13663_),
    .A3(_13672_),
    .A4(_13683_),
    .ZN(_13684_));
 OR2_X2 _23379_ (.A1(_13684_),
    .A2(_11775_),
    .ZN(_13685_));
 XOR2_X2 _23380_ (.A(_13637_),
    .B(_13685_),
    .Z(_13686_));
 AOI21_X1 _23381_ (.A(_13053_),
    .B1(_11441_),
    .B2(_11328_),
    .ZN(_13687_));
 AOI21_X1 _23382_ (.A(_13687_),
    .B1(_11540_),
    .B2(_12374_),
    .ZN(_13688_));
 OAI21_X1 _23383_ (.A(_12374_),
    .B1(_12375_),
    .B2(_11425_),
    .ZN(_13689_));
 OAI21_X1 _23384_ (.A(_12374_),
    .B1(_12338_),
    .B2(_12322_),
    .ZN(_13690_));
 AND3_X1 _23385_ (.A1(_13688_),
    .A2(_13689_),
    .A3(_13690_),
    .ZN(_13691_));
 OAI21_X1 _23386_ (.A(_11415_),
    .B1(_11444_),
    .B2(_12324_),
    .ZN(_13692_));
 OAI21_X1 _23387_ (.A(_11415_),
    .B1(_12375_),
    .B2(_13070_),
    .ZN(_13693_));
 INV_X1 _23388_ (.A(_12720_),
    .ZN(_13694_));
 NOR4_X1 _23389_ (.A1(_13694_),
    .A2(_13078_),
    .A3(_11449_),
    .A4(_13080_),
    .ZN(_13695_));
 AND4_X1 _23390_ (.A1(_13691_),
    .A2(_13692_),
    .A3(_13693_),
    .A4(_13695_),
    .ZN(_13696_));
 NAND3_X1 _23391_ (.A1(_12369_),
    .A2(_12666_),
    .A3(_13067_),
    .ZN(_13697_));
 AND2_X1 _23392_ (.A1(_11533_),
    .A2(_11369_),
    .ZN(_13698_));
 OR3_X1 _23393_ (.A1(_13527_),
    .A2(_13698_),
    .A3(_13529_),
    .ZN(_13699_));
 NOR3_X1 _23394_ (.A1(_13697_),
    .A2(_13699_),
    .A3(_12355_),
    .ZN(_13700_));
 OAI22_X1 _23395_ (.A1(_11440_),
    .A2(_11341_),
    .B1(_12297_),
    .B2(_12697_),
    .ZN(_13701_));
 AND2_X1 _23396_ (.A1(_11331_),
    .A2(_11425_),
    .ZN(_13702_));
 AND2_X1 _23397_ (.A1(_11467_),
    .A2(_11405_),
    .ZN(_13703_));
 OR4_X1 _23398_ (.A1(_13549_),
    .A2(_13701_),
    .A3(_13702_),
    .A4(_13703_),
    .ZN(_13704_));
 OAI21_X1 _23399_ (.A(_11353_),
    .B1(_12324_),
    .B2(_13070_),
    .ZN(_13705_));
 NAND3_X1 _23400_ (.A1(_13340_),
    .A2(_13315_),
    .A3(_13705_),
    .ZN(_13706_));
 NOR4_X1 _23401_ (.A1(_13704_),
    .A2(_11348_),
    .A3(_11339_),
    .A4(_13706_),
    .ZN(_13707_));
 NAND2_X1 _23402_ (.A1(_11540_),
    .A2(_11497_),
    .ZN(_13708_));
 NAND2_X1 _23403_ (.A1(_11386_),
    .A2(_11530_),
    .ZN(_13709_));
 NAND3_X1 _23404_ (.A1(_13708_),
    .A2(_13709_),
    .A3(_11516_),
    .ZN(_13710_));
 OAI22_X1 _23405_ (.A1(_12715_),
    .A2(_12329_),
    .B1(_12694_),
    .B2(_12318_),
    .ZN(_13711_));
 NOR4_X1 _23406_ (.A1(_13710_),
    .A2(_11438_),
    .A3(_12654_),
    .A4(_13711_),
    .ZN(_13712_));
 NAND4_X1 _23407_ (.A1(_13696_),
    .A2(_13700_),
    .A3(_13707_),
    .A4(_13712_),
    .ZN(_13713_));
 AND3_X1 _23408_ (.A1(_11534_),
    .A2(_12324_),
    .A3(_11338_),
    .ZN(_13714_));
 OAI21_X1 _23409_ (.A(_13316_),
    .B1(_12297_),
    .B2(_12287_),
    .ZN(_13715_));
 AOI211_X1 _23410_ (.A(_13714_),
    .B(_13715_),
    .C1(_11472_),
    .C2(_11514_),
    .ZN(_13716_));
 NOR3_X1 _23411_ (.A1(_11495_),
    .A2(_12363_),
    .A3(_11428_),
    .ZN(_13717_));
 AOI22_X1 _23412_ (.A1(_11482_),
    .A2(_12322_),
    .B1(_11370_),
    .B2(_11483_),
    .ZN(_13718_));
 AOI22_X1 _23413_ (.A1(_11493_),
    .A2(_11482_),
    .B1(_12375_),
    .B2(_11497_),
    .ZN(_13719_));
 AND4_X1 _23414_ (.A1(_13716_),
    .A2(_13717_),
    .A3(_13718_),
    .A4(_13719_),
    .ZN(_13720_));
 AOI221_X4 _23415_ (.A(_13556_),
    .B1(_11536_),
    .B2(_11452_),
    .C1(_11540_),
    .C2(_11460_),
    .ZN(_13721_));
 OR2_X1 _23416_ (.A1(_12313_),
    .A2(_11447_),
    .ZN(_13722_));
 NAND2_X1 _23417_ (.A1(_12366_),
    .A2(_11525_),
    .ZN(_13723_));
 OAI21_X1 _23418_ (.A(_13723_),
    .B1(_12345_),
    .B2(_11328_),
    .ZN(_13724_));
 AND2_X1 _23419_ (.A1(_11481_),
    .A2(_11371_),
    .ZN(_13725_));
 AND2_X1 _23420_ (.A1(_11450_),
    .A2(_13070_),
    .ZN(_13726_));
 NOR4_X1 _23421_ (.A1(_13724_),
    .A2(_13725_),
    .A3(_13550_),
    .A4(_13726_),
    .ZN(_13727_));
 OAI21_X1 _23422_ (.A(_11431_),
    .B1(_11493_),
    .B2(_11467_),
    .ZN(_13728_));
 NAND3_X1 _23423_ (.A1(_11353_),
    .A2(_13036_),
    .A3(_12690_),
    .ZN(_13729_));
 AND4_X1 _23424_ (.A1(_13722_),
    .A2(_13727_),
    .A3(_13728_),
    .A4(_13729_),
    .ZN(_13730_));
 NAND2_X1 _23425_ (.A1(_11406_),
    .A2(_11393_),
    .ZN(_13731_));
 OAI21_X1 _23426_ (.A(_11460_),
    .B1(_11344_),
    .B2(_12375_),
    .ZN(_13732_));
 AOI22_X1 _23427_ (.A1(_12338_),
    .A2(_11431_),
    .B1(_11403_),
    .B2(_11528_),
    .ZN(_13733_));
 AND4_X1 _23428_ (.A1(_13731_),
    .A2(_13049_),
    .A3(_13732_),
    .A4(_13733_),
    .ZN(_13734_));
 NAND4_X1 _23429_ (.A1(_13720_),
    .A2(_13721_),
    .A3(_13730_),
    .A4(_13734_),
    .ZN(_13735_));
 NOR2_X2 _23430_ (.A1(_13713_),
    .A2(_13735_),
    .ZN(_13736_));
 XNOR2_X1 _23431_ (.A(_13463_),
    .B(_13736_),
    .ZN(_13737_));
 XNOR2_X1 _23432_ (.A(_13686_),
    .B(_13737_),
    .ZN(_13738_));
 NOR2_X1 _23433_ (.A1(_12443_),
    .A2(_13484_),
    .ZN(_13739_));
 NAND2_X1 _23434_ (.A1(_12417_),
    .A2(_12391_),
    .ZN(_13740_));
 AND4_X1 _23435_ (.A1(_12005_),
    .A2(_13739_),
    .A3(_13740_),
    .A4(_12393_),
    .ZN(_13741_));
 OAI21_X1 _23436_ (.A(_12078_),
    .B1(_11894_),
    .B2(_12449_),
    .ZN(_13742_));
 NAND2_X1 _23437_ (.A1(_12795_),
    .A2(_13742_),
    .ZN(_13743_));
 OR4_X1 _23438_ (.A1(_12460_),
    .A2(_13743_),
    .A3(_12759_),
    .A4(_12757_),
    .ZN(_13744_));
 AOI22_X1 _23439_ (.A1(_12737_),
    .A2(_12009_),
    .B1(_11983_),
    .B2(_11985_),
    .ZN(_13745_));
 OAI221_X1 _23440_ (.A(_13745_),
    .B1(_12387_),
    .B2(_12740_),
    .C1(_12388_),
    .C2(_12458_),
    .ZN(_13746_));
 AOI21_X1 _23441_ (.A(_12753_),
    .B1(_12400_),
    .B2(_13271_),
    .ZN(_13747_));
 NOR4_X1 _23442_ (.A1(_13744_),
    .A2(_13746_),
    .A3(_12995_),
    .A4(_13747_),
    .ZN(_13748_));
 AND2_X1 _23443_ (.A1(_11974_),
    .A2(_11987_),
    .ZN(_13749_));
 INV_X1 _23444_ (.A(_13749_),
    .ZN(_13750_));
 OAI211_X1 _23445_ (.A(_13750_),
    .B(_13473_),
    .C1(_11935_),
    .C2(_12039_),
    .ZN(_13751_));
 AOI22_X1 _23446_ (.A1(_12762_),
    .A2(_12034_),
    .B1(_12763_),
    .B2(_11926_),
    .ZN(_13752_));
 NAND2_X1 _23447_ (.A1(_11964_),
    .A2(_12088_),
    .ZN(_13753_));
 OAI211_X1 _23448_ (.A(_13752_),
    .B(_13753_),
    .C1(_12045_),
    .C2(_12742_),
    .ZN(_13754_));
 AND3_X1 _23449_ (.A1(_12391_),
    .A2(_11906_),
    .A3(_12011_),
    .ZN(_13755_));
 OAI21_X1 _23450_ (.A(_12009_),
    .B1(_12763_),
    .B2(_11987_),
    .ZN(_13756_));
 OAI211_X1 _23451_ (.A(_13756_),
    .B(_13489_),
    .C1(_12039_),
    .C2(_12458_),
    .ZN(_13757_));
 NOR4_X1 _23452_ (.A1(_13751_),
    .A2(_13754_),
    .A3(_13755_),
    .A4(_13757_),
    .ZN(_13758_));
 OAI21_X1 _23453_ (.A(_12094_),
    .B1(_11930_),
    .B2(_12010_),
    .ZN(_13759_));
 AOI21_X1 _23454_ (.A(_12069_),
    .B1(_12083_),
    .B2(_12388_),
    .ZN(_13760_));
 OAI21_X1 _23455_ (.A(_12074_),
    .B1(_12069_),
    .B2(_11938_),
    .ZN(_13761_));
 NOR4_X1 _23456_ (.A1(_13760_),
    .A2(_13761_),
    .A3(_13283_),
    .A4(_12498_),
    .ZN(_13762_));
 OAI21_X1 _23457_ (.A(_11993_),
    .B1(_11929_),
    .B2(_12090_),
    .ZN(_13763_));
 OAI211_X1 _23458_ (.A(_11941_),
    .B(_11979_),
    .C1(_11980_),
    .C2(_12410_),
    .ZN(_13764_));
 AND4_X1 _23459_ (.A1(_13759_),
    .A2(_13762_),
    .A3(_13763_),
    .A4(_13764_),
    .ZN(_13765_));
 AND4_X1 _23460_ (.A1(_13741_),
    .A2(_13748_),
    .A3(_13758_),
    .A4(_13765_),
    .ZN(_13766_));
 AOI21_X1 _23461_ (.A(_12475_),
    .B1(_12743_),
    .B2(_12387_),
    .ZN(_13767_));
 NAND2_X1 _23462_ (.A1(_12009_),
    .A2(_12412_),
    .ZN(_13768_));
 NAND2_X1 _23463_ (.A1(_12461_),
    .A2(_12024_),
    .ZN(_13769_));
 NAND2_X1 _23464_ (.A1(_13768_),
    .A2(_13769_),
    .ZN(_13770_));
 NOR3_X1 _23465_ (.A1(_12436_),
    .A2(_13767_),
    .A3(_13770_),
    .ZN(_13771_));
 OAI221_X1 _23466_ (.A(_11976_),
    .B1(_12432_),
    .B2(_12753_),
    .C1(_12406_),
    .C2(_12445_),
    .ZN(_13772_));
 INV_X1 _23467_ (.A(_13466_),
    .ZN(_13773_));
 OAI21_X1 _23468_ (.A(_13773_),
    .B1(_12044_),
    .B2(_12395_),
    .ZN(_13774_));
 AND2_X1 _23469_ (.A1(_12064_),
    .A2(_12084_),
    .ZN(_13775_));
 NAND3_X1 _23470_ (.A1(_12739_),
    .A2(_13498_),
    .A3(_13509_),
    .ZN(_13776_));
 NOR4_X1 _23471_ (.A1(_13772_),
    .A2(_13774_),
    .A3(_13775_),
    .A4(_13776_),
    .ZN(_13777_));
 OAI21_X1 _23472_ (.A(_12489_),
    .B1(_11937_),
    .B2(_11930_),
    .ZN(_13778_));
 AOI221_X4 _23473_ (.A(_11901_),
    .B1(_11959_),
    .B2(_11950_),
    .C1(_12024_),
    .C2(_12088_),
    .ZN(_13779_));
 AOI22_X1 _23474_ (.A1(_11959_),
    .A2(_12737_),
    .B1(_11952_),
    .B2(_11942_),
    .ZN(_13780_));
 NAND2_X1 _23475_ (.A1(_12080_),
    .A2(_11926_),
    .ZN(_13781_));
 AND3_X1 _23476_ (.A1(_13780_),
    .A2(_11965_),
    .A3(_13781_),
    .ZN(_13782_));
 AND4_X1 _23477_ (.A1(_13778_),
    .A2(_13779_),
    .A3(_12021_),
    .A4(_13782_),
    .ZN(_13783_));
 AOI22_X1 _23478_ (.A1(_11974_),
    .A2(_11937_),
    .B1(_12480_),
    .B2(_12401_),
    .ZN(_13784_));
 OAI211_X1 _23479_ (.A(_13784_),
    .B(_13273_),
    .C1(_12402_),
    .C2(_12753_),
    .ZN(_13785_));
 AND2_X1 _23480_ (.A1(_11980_),
    .A2(_12030_),
    .ZN(_13786_));
 OR2_X1 _23481_ (.A1(_12031_),
    .A2(_13786_),
    .ZN(_13787_));
 OAI211_X1 _23482_ (.A(_12444_),
    .B(_12053_),
    .C1(_12044_),
    .C2(_12388_),
    .ZN(_13788_));
 NOR4_X1 _23483_ (.A1(_13785_),
    .A2(_12042_),
    .A3(_13787_),
    .A4(_13788_),
    .ZN(_13789_));
 AND4_X1 _23484_ (.A1(_13771_),
    .A2(_13777_),
    .A3(_13783_),
    .A4(_13789_),
    .ZN(_13790_));
 NAND2_X2 _23485_ (.A1(_13766_),
    .A2(_13790_),
    .ZN(_13791_));
 XNOR2_X1 _23486_ (.A(_13738_),
    .B(_13791_),
    .ZN(_13792_));
 INV_X1 _23487_ (.A(_17191_),
    .ZN(_13793_));
 XNOR2_X1 _23488_ (.A(_13792_),
    .B(_13793_),
    .ZN(_13794_));
 MUX2_X1 _23489_ (.A(_13584_),
    .B(_13794_),
    .S(_11084_),
    .Z(_00722_));
 XOR2_X1 _23490_ (.A(_17192_),
    .B(_16995_),
    .Z(_13795_));
 OAI21_X1 _23491_ (.A(_11460_),
    .B1(_11489_),
    .B2(_13084_),
    .ZN(_13796_));
 AOI21_X1 _23492_ (.A(_11440_),
    .B1(_11539_),
    .B2(_12715_),
    .ZN(_13797_));
 AOI211_X1 _23493_ (.A(_13550_),
    .B(_13797_),
    .C1(_11420_),
    .C2(_11366_),
    .ZN(_13798_));
 OAI21_X1 _23494_ (.A(_11460_),
    .B1(_11437_),
    .B2(_11505_),
    .ZN(_13799_));
 NOR2_X1 _23495_ (.A1(_12302_),
    .A2(_11367_),
    .ZN(_13800_));
 AND4_X1 _23496_ (.A1(_13796_),
    .A2(_13798_),
    .A3(_13799_),
    .A4(_13800_),
    .ZN(_13801_));
 NAND2_X1 _23497_ (.A1(_11431_),
    .A2(_11442_),
    .ZN(_13802_));
 OAI21_X1 _23498_ (.A(_11414_),
    .B1(_11370_),
    .B2(_11371_),
    .ZN(_13803_));
 AND4_X1 _23499_ (.A1(_13332_),
    .A2(_13334_),
    .A3(_13034_),
    .A4(_13803_),
    .ZN(_13804_));
 AOI211_X1 _23500_ (.A(_11474_),
    .B(_11430_),
    .C1(_12337_),
    .C2(_11427_),
    .ZN(_13805_));
 AND4_X1 _23501_ (.A1(_13802_),
    .A2(_13804_),
    .A3(_13805_),
    .A4(_12701_),
    .ZN(_13806_));
 AND3_X1 _23502_ (.A1(_11521_),
    .A2(_13036_),
    .A3(_12664_),
    .ZN(_13807_));
 AOI21_X1 _23503_ (.A(_13807_),
    .B1(_11522_),
    .B2(_12717_),
    .ZN(_13808_));
 OAI21_X1 _23504_ (.A(_11522_),
    .B1(_11518_),
    .B2(_11530_),
    .ZN(_13809_));
 OAI21_X1 _23505_ (.A(_11353_),
    .B1(_11444_),
    .B2(_11400_),
    .ZN(_13810_));
 AND4_X1 _23506_ (.A1(_12704_),
    .A2(_13808_),
    .A3(_13809_),
    .A4(_13810_),
    .ZN(_13811_));
 AND3_X1 _23507_ (.A1(_11477_),
    .A2(_11408_),
    .A3(_11423_),
    .ZN(_13812_));
 OR4_X1 _23508_ (.A1(_12368_),
    .A2(_13812_),
    .A3(_12667_),
    .A4(_13527_),
    .ZN(_13813_));
 OR2_X1 _23509_ (.A1(_12652_),
    .A2(_13528_),
    .ZN(_13814_));
 AND2_X1 _23510_ (.A1(_11382_),
    .A2(_11327_),
    .ZN(_13815_));
 NOR4_X1 _23511_ (.A1(_13813_),
    .A2(_11383_),
    .A3(_13814_),
    .A4(_13815_),
    .ZN(_13816_));
 NAND4_X2 _23512_ (.A1(_13801_),
    .A2(_13806_),
    .A3(_13811_),
    .A4(_13816_),
    .ZN(_13817_));
 AOI211_X1 _23513_ (.A(_11378_),
    .B(_12697_),
    .C1(_11338_),
    .C2(_11360_),
    .ZN(_13818_));
 NOR4_X1 _23514_ (.A1(_13818_),
    .A2(_13296_),
    .A3(_12355_),
    .A4(_11531_),
    .ZN(_13819_));
 OAI211_X1 _23515_ (.A(_11317_),
    .B(_11395_),
    .C1(_11418_),
    .C2(_11361_),
    .ZN(_13820_));
 NAND4_X1 _23516_ (.A1(_11314_),
    .A2(_11316_),
    .A3(_11335_),
    .A4(_11320_),
    .ZN(_13821_));
 AND2_X1 _23517_ (.A1(_13820_),
    .A2(_13821_),
    .ZN(_13822_));
 OAI21_X1 _23518_ (.A(_11318_),
    .B1(_12717_),
    .B2(_11369_),
    .ZN(_13823_));
 OAI21_X1 _23519_ (.A(_11450_),
    .B1(_11492_),
    .B2(_11467_),
    .ZN(_13824_));
 OAI21_X1 _23520_ (.A(_11450_),
    .B1(_12321_),
    .B2(_11456_),
    .ZN(_13825_));
 AND4_X1 _23521_ (.A1(_13822_),
    .A2(_13823_),
    .A3(_13824_),
    .A4(_13825_),
    .ZN(_13826_));
 OAI21_X1 _23522_ (.A(_11331_),
    .B1(_11467_),
    .B2(_11389_),
    .ZN(_13827_));
 OAI21_X1 _23523_ (.A(_11331_),
    .B1(_11489_),
    .B2(_11525_),
    .ZN(_13828_));
 AND4_X1 _23524_ (.A1(_13819_),
    .A2(_13826_),
    .A3(_13827_),
    .A4(_13828_),
    .ZN(_13829_));
 NAND3_X1 _23525_ (.A1(_11380_),
    .A2(_13036_),
    .A3(_11488_),
    .ZN(_13830_));
 AND2_X1 _23526_ (.A1(_11419_),
    .A2(_11533_),
    .ZN(_13831_));
 AOI211_X1 _23527_ (.A(_13831_),
    .B(_13548_),
    .C1(_11534_),
    .C2(_11327_),
    .ZN(_13832_));
 OAI211_X1 _23528_ (.A(_11487_),
    .B(_11423_),
    .C1(_11435_),
    .C2(_11472_),
    .ZN(_13833_));
 AND2_X1 _23529_ (.A1(_11533_),
    .A2(_12321_),
    .ZN(_13834_));
 AND2_X1 _23530_ (.A1(_12337_),
    .A2(_11533_),
    .ZN(_13835_));
 NOR4_X1 _23531_ (.A1(_13834_),
    .A2(_13835_),
    .A3(_12659_),
    .A4(_13698_),
    .ZN(_13836_));
 AND4_X1 _23532_ (.A1(_13830_),
    .A2(_13832_),
    .A3(_13833_),
    .A4(_13836_),
    .ZN(_13837_));
 NOR4_X1 _23533_ (.A1(_11508_),
    .A2(_12713_),
    .A3(_13087_),
    .A4(_11506_),
    .ZN(_13838_));
 OAI21_X1 _23534_ (.A(_11386_),
    .B1(_12322_),
    .B2(_13084_),
    .ZN(_13839_));
 AND3_X1 _23535_ (.A1(_13839_),
    .A2(_13709_),
    .A3(_12331_),
    .ZN(_13840_));
 NAND4_X2 _23536_ (.A1(_13829_),
    .A2(_13837_),
    .A3(_13838_),
    .A4(_13840_),
    .ZN(_13841_));
 NOR2_X4 _23537_ (.A1(_13817_),
    .A2(_13841_),
    .ZN(_13842_));
 XNOR2_X1 _23538_ (.A(_13685_),
    .B(_13842_),
    .ZN(_13843_));
 NAND3_X1 _23539_ (.A1(_12226_),
    .A2(_11255_),
    .A3(_11091_),
    .ZN(_13844_));
 AND3_X1 _23540_ (.A1(_11103_),
    .A2(_11099_),
    .A3(_11270_),
    .ZN(_13845_));
 NOR4_X1 _23541_ (.A1(_13189_),
    .A2(_12234_),
    .A3(_12235_),
    .A4(_13845_),
    .ZN(_13846_));
 OAI211_X1 _23542_ (.A(_11255_),
    .B(_11091_),
    .C1(_11181_),
    .C2(_11160_),
    .ZN(_13847_));
 OAI21_X1 _23543_ (.A(_11092_),
    .B1(_12829_),
    .B2(_11235_),
    .ZN(_13848_));
 AND4_X1 _23544_ (.A1(_13844_),
    .A2(_13846_),
    .A3(_13847_),
    .A4(_13848_),
    .ZN(_13849_));
 AOI21_X1 _23545_ (.A(_12224_),
    .B1(_12260_),
    .B2(_11178_),
    .ZN(_13850_));
 AOI21_X1 _23546_ (.A(_13850_),
    .B1(_11149_),
    .B2(_11096_),
    .ZN(_13851_));
 OAI21_X1 _23547_ (.A(_11148_),
    .B1(_12580_),
    .B2(_11163_),
    .ZN(_13852_));
 OAI21_X1 _23548_ (.A(_11136_),
    .B1(_12275_),
    .B2(_12226_),
    .ZN(_13853_));
 OAI21_X1 _23549_ (.A(_11136_),
    .B1(_11304_),
    .B2(_11286_),
    .ZN(_13854_));
 AND4_X1 _23550_ (.A1(_13851_),
    .A2(_13852_),
    .A3(_13853_),
    .A4(_13854_),
    .ZN(_13855_));
 NAND4_X1 _23551_ (.A1(_12182_),
    .A2(_11155_),
    .A3(_11170_),
    .A4(_11153_),
    .ZN(_13856_));
 OAI211_X1 _23552_ (.A(_13369_),
    .B(_13856_),
    .C1(_11209_),
    .C2(_11111_),
    .ZN(_13857_));
 AND4_X1 _23553_ (.A1(_11203_),
    .A2(_11171_),
    .A3(_11098_),
    .A4(_11270_),
    .ZN(_13858_));
 AND3_X1 _23554_ (.A1(_11171_),
    .A2(_11126_),
    .A3(_11118_),
    .ZN(_13859_));
 OR3_X1 _23555_ (.A1(_13858_),
    .A2(_13859_),
    .A3(_12247_),
    .ZN(_13860_));
 OAI21_X1 _23556_ (.A(_12242_),
    .B1(_12251_),
    .B2(_11209_),
    .ZN(_13861_));
 AOI21_X1 _23557_ (.A(_11209_),
    .B1(_12229_),
    .B2(_11293_),
    .ZN(_13862_));
 NOR4_X1 _23558_ (.A1(_13857_),
    .A2(_13860_),
    .A3(_13861_),
    .A4(_13862_),
    .ZN(_13863_));
 OAI21_X1 _23559_ (.A(_11199_),
    .B1(_11304_),
    .B2(_12830_),
    .ZN(_13864_));
 OAI21_X1 _23560_ (.A(_11213_),
    .B1(_11225_),
    .B2(_11128_),
    .ZN(_13865_));
 OAI21_X1 _23561_ (.A(_11213_),
    .B1(_11152_),
    .B2(_11223_),
    .ZN(_13866_));
 OAI211_X1 _23562_ (.A(_11199_),
    .B(_11095_),
    .C1(_11153_),
    .C2(_11099_),
    .ZN(_13867_));
 AND4_X1 _23563_ (.A1(_13864_),
    .A2(_13865_),
    .A3(_13866_),
    .A4(_13867_),
    .ZN(_13868_));
 NAND4_X2 _23564_ (.A1(_13849_),
    .A2(_13855_),
    .A3(_13863_),
    .A4(_13868_),
    .ZN(_13869_));
 OAI21_X1 _23565_ (.A(_13390_),
    .B1(_11276_),
    .B2(_11268_),
    .ZN(_13870_));
 NOR3_X1 _23566_ (.A1(_11189_),
    .A2(_11097_),
    .A3(_16738_),
    .ZN(_13871_));
 AND3_X1 _23567_ (.A1(_13871_),
    .A2(_11088_),
    .A3(_11263_),
    .ZN(_13872_));
 NOR4_X1 _23568_ (.A1(_13870_),
    .A2(_12200_),
    .A3(_11275_),
    .A4(_13872_),
    .ZN(_13873_));
 OAI21_X1 _23569_ (.A(_11297_),
    .B1(_11282_),
    .B2(_11223_),
    .ZN(_13874_));
 AND4_X1 _23570_ (.A1(_12857_),
    .A2(_13873_),
    .A3(_13393_),
    .A4(_13874_),
    .ZN(_13875_));
 AND2_X1 _23571_ (.A1(_13173_),
    .A2(_13174_),
    .ZN(_13876_));
 AND2_X1 _23572_ (.A1(_11127_),
    .A2(_11291_),
    .ZN(_13877_));
 AOI211_X1 _23573_ (.A(_12196_),
    .B(_13877_),
    .C1(_11302_),
    .C2(_11291_),
    .ZN(_13878_));
 OAI21_X1 _23574_ (.A(_11291_),
    .B1(_13871_),
    .B2(_11248_),
    .ZN(_13879_));
 OAI21_X1 _23575_ (.A(_11264_),
    .B1(_12199_),
    .B2(_11116_),
    .ZN(_13880_));
 AND4_X1 _23576_ (.A1(_13876_),
    .A2(_13878_),
    .A3(_13879_),
    .A4(_13880_),
    .ZN(_13881_));
 OAI21_X1 _23577_ (.A(_11252_),
    .B1(_12580_),
    .B2(_12230_),
    .ZN(_13882_));
 OAI21_X1 _23578_ (.A(_11252_),
    .B1(_11152_),
    .B2(_11096_),
    .ZN(_13883_));
 OAI21_X1 _23579_ (.A(_11234_),
    .B1(_11279_),
    .B2(_11177_),
    .ZN(_13884_));
 AND4_X1 _23580_ (.A1(_12609_),
    .A2(_13882_),
    .A3(_13883_),
    .A4(_13884_),
    .ZN(_13885_));
 OAI211_X1 _23581_ (.A(_11088_),
    .B(_11237_),
    .C1(_11301_),
    .C2(_12187_),
    .ZN(_13886_));
 OAI211_X1 _23582_ (.A(_11088_),
    .B(_11237_),
    .C1(_11121_),
    .C2(_11139_),
    .ZN(_13887_));
 OAI211_X1 _23583_ (.A(_13886_),
    .B(_13887_),
    .C1(_12588_),
    .C2(_11278_),
    .ZN(_13888_));
 NAND3_X1 _23584_ (.A1(_11121_),
    .A2(_11237_),
    .A3(_11102_),
    .ZN(_13889_));
 NAND3_X1 _23585_ (.A1(_11304_),
    .A2(_11237_),
    .A3(_11102_),
    .ZN(_13890_));
 NAND2_X1 _23586_ (.A1(_13889_),
    .A2(_13890_),
    .ZN(_13891_));
 AND2_X1 _23587_ (.A1(_11243_),
    .A2(_11160_),
    .ZN(_13892_));
 NOR4_X1 _23588_ (.A1(_13888_),
    .A2(_13891_),
    .A3(_11244_),
    .A4(_13892_),
    .ZN(_13893_));
 NAND4_X2 _23589_ (.A1(_13875_),
    .A2(_13881_),
    .A3(_13885_),
    .A4(_13893_),
    .ZN(_13894_));
 NOR2_X4 _23590_ (.A1(_13869_),
    .A2(_13894_),
    .ZN(_13895_));
 XOR2_X2 _23591_ (.A(_13895_),
    .B(_11877_),
    .Z(_13896_));
 XNOR2_X1 _23592_ (.A(_13843_),
    .B(_13896_),
    .ZN(_13897_));
 AND3_X1 _23593_ (.A1(_12730_),
    .A2(_12026_),
    .A3(_13486_),
    .ZN(_13898_));
 OAI21_X1 _23594_ (.A(_12022_),
    .B1(_12401_),
    .B2(_12455_),
    .ZN(_13899_));
 OAI211_X1 _23595_ (.A(_13898_),
    .B(_13899_),
    .C1(_12013_),
    .C2(_12044_),
    .ZN(_13900_));
 AND2_X1 _23596_ (.A1(_12088_),
    .A2(_12058_),
    .ZN(_13901_));
 OAI211_X1 _23597_ (.A(_13753_),
    .B(_13266_),
    .C1(_12071_),
    .C2(_12742_),
    .ZN(_13902_));
 AOI21_X1 _23598_ (.A(_12756_),
    .B1(_12081_),
    .B2(_12406_),
    .ZN(_13903_));
 AOI21_X1 _23599_ (.A(_12756_),
    .B1(_12083_),
    .B2(_12036_),
    .ZN(_13904_));
 OR4_X1 _23600_ (.A1(_13901_),
    .A2(_13902_),
    .A3(_13903_),
    .A4(_13904_),
    .ZN(_13905_));
 NOR2_X1 _23601_ (.A1(_12037_),
    .A2(_12496_),
    .ZN(_13906_));
 NOR4_X1 _23602_ (.A1(_13900_),
    .A2(_13905_),
    .A3(_13906_),
    .A4(_13012_),
    .ZN(_13907_));
 AND2_X1 _23603_ (.A1(_12801_),
    .A2(_12429_),
    .ZN(_13908_));
 OR4_X1 _23604_ (.A1(_12776_),
    .A2(_13908_),
    .A3(_12960_),
    .A4(_13749_),
    .ZN(_13909_));
 OAI21_X1 _23605_ (.A(_11993_),
    .B1(_11989_),
    .B2(_12780_),
    .ZN(_13910_));
 OAI211_X1 _23606_ (.A(_11941_),
    .B(_11979_),
    .C1(_11980_),
    .C2(_12024_),
    .ZN(_13911_));
 OAI211_X1 _23607_ (.A(_13910_),
    .B(_13911_),
    .C1(_11984_),
    .C2(_13271_),
    .ZN(_13912_));
 NAND4_X1 _23608_ (.A1(_13237_),
    .A2(_12008_),
    .A3(_13768_),
    .A4(_12803_),
    .ZN(_13913_));
 OAI21_X1 _23609_ (.A(_12461_),
    .B1(_12737_),
    .B2(_11898_),
    .ZN(_13914_));
 OAI21_X1 _23610_ (.A(_12461_),
    .B1(_12090_),
    .B2(_11994_),
    .ZN(_13915_));
 OAI211_X1 _23611_ (.A(_11924_),
    .B(_11979_),
    .C1(_12447_),
    .C2(_11900_),
    .ZN(_13916_));
 NAND4_X1 _23612_ (.A1(_13914_),
    .A2(_13915_),
    .A3(_13769_),
    .A4(_13916_),
    .ZN(_13917_));
 NOR4_X1 _23613_ (.A1(_13909_),
    .A2(_13912_),
    .A3(_13913_),
    .A4(_13917_),
    .ZN(_13918_));
 NAND2_X1 _23614_ (.A1(_11952_),
    .A2(_12078_),
    .ZN(_13919_));
 OAI21_X1 _23615_ (.A(_13919_),
    .B1(_12079_),
    .B2(_13271_),
    .ZN(_13920_));
 AOI21_X1 _23616_ (.A(_13920_),
    .B1(_12078_),
    .B2(_12399_),
    .ZN(_13921_));
 AND3_X1 _23617_ (.A1(_12068_),
    .A2(_11955_),
    .A3(_12429_),
    .ZN(_13922_));
 NOR4_X1 _23618_ (.A1(_13281_),
    .A2(_13922_),
    .A3(_12783_),
    .A4(_13284_),
    .ZN(_13923_));
 OAI21_X1 _23619_ (.A(_12064_),
    .B1(_12438_),
    .B2(_12410_),
    .ZN(_13924_));
 NAND2_X1 _23620_ (.A1(_12064_),
    .A2(_11937_),
    .ZN(_13925_));
 OAI21_X1 _23621_ (.A(_12064_),
    .B1(_12447_),
    .B2(_11900_),
    .ZN(_13926_));
 AND3_X1 _23622_ (.A1(_13924_),
    .A2(_13925_),
    .A3(_13926_),
    .ZN(_13927_));
 NAND2_X1 _23623_ (.A1(_12033_),
    .A2(_12440_),
    .ZN(_13928_));
 AND4_X1 _23624_ (.A1(_13928_),
    .A2(_12052_),
    .A3(_12056_),
    .A4(_13477_),
    .ZN(_13929_));
 AND4_X1 _23625_ (.A1(_13921_),
    .A2(_13923_),
    .A3(_13927_),
    .A4(_13929_),
    .ZN(_13930_));
 INV_X1 _23626_ (.A(_12954_),
    .ZN(_13931_));
 AND2_X1 _23627_ (.A1(_11964_),
    .A2(_11887_),
    .ZN(_13932_));
 OR4_X1 _23628_ (.A1(_13931_),
    .A2(_11901_),
    .A3(_13932_),
    .A4(_12478_),
    .ZN(_13933_));
 OAI21_X1 _23629_ (.A(_12480_),
    .B1(_11953_),
    .B2(_13270_),
    .ZN(_13934_));
 OAI211_X1 _23630_ (.A(_11977_),
    .B(_11912_),
    .C1(_12447_),
    .C2(_11987_),
    .ZN(_13935_));
 NAND4_X1 _23631_ (.A1(_11977_),
    .A2(_12414_),
    .A3(_11932_),
    .A4(_11912_),
    .ZN(_13936_));
 NAND3_X1 _23632_ (.A1(_13934_),
    .A2(_13935_),
    .A3(_13936_),
    .ZN(_13937_));
 INV_X1 _23633_ (.A(_11951_),
    .ZN(_13938_));
 OAI21_X1 _23634_ (.A(_11943_),
    .B1(_12033_),
    .B2(_12080_),
    .ZN(_13939_));
 NAND4_X1 _23635_ (.A1(_13938_),
    .A2(_12752_),
    .A3(_12972_),
    .A4(_13939_),
    .ZN(_13940_));
 OAI21_X1 _23636_ (.A(_12489_),
    .B1(_11953_),
    .B2(_12027_),
    .ZN(_13941_));
 OAI211_X1 _23637_ (.A(_12489_),
    .B(_11944_),
    .C1(_11919_),
    .C2(_11920_),
    .ZN(_13942_));
 OAI211_X1 _23638_ (.A(_13941_),
    .B(_13942_),
    .C1(_11935_),
    .C2(_11991_),
    .ZN(_13943_));
 NOR4_X1 _23639_ (.A1(_13933_),
    .A2(_13937_),
    .A3(_13940_),
    .A4(_13943_),
    .ZN(_13944_));
 AND4_X1 _23640_ (.A1(_13907_),
    .A2(_13918_),
    .A3(_13930_),
    .A4(_13944_),
    .ZN(_13945_));
 NAND2_X2 _23641_ (.A1(_13945_),
    .A2(_12778_),
    .ZN(_13946_));
 XNOR2_X1 _23642_ (.A(_13897_),
    .B(_13946_),
    .ZN(_13947_));
 XOR2_X1 _23643_ (.A(_13947_),
    .B(_17192_),
    .Z(_13948_));
 MUX2_X1 _23644_ (.A(_13795_),
    .B(_13948_),
    .S(_11084_),
    .Z(_00723_));
 AND2_X2 _23645_ (.A1(_17087_),
    .A2(_17088_),
    .ZN(_13949_));
 AND2_X1 _23646_ (.A1(_17090_),
    .A2(_17091_),
    .ZN(_13950_));
 AND2_X1 _23647_ (.A1(_13949_),
    .A2(_13950_),
    .ZN(_13951_));
 BUF_X2 _23648_ (.A(_13951_),
    .Z(_13952_));
 BUF_X2 _23649_ (.A(_13952_),
    .Z(_13953_));
 INV_X1 _23650_ (.A(_17084_),
    .ZN(_13954_));
 NOR2_X2 _23651_ (.A1(_13954_),
    .A2(_17083_),
    .ZN(_13955_));
 AND2_X1 _23652_ (.A1(_17085_),
    .A2(_17086_),
    .ZN(_13956_));
 CLKBUF_X2 _23653_ (.A(_13956_),
    .Z(_13957_));
 AND2_X1 _23654_ (.A1(_13955_),
    .A2(_13957_),
    .ZN(_13958_));
 BUF_X2 _23655_ (.A(_13958_),
    .Z(_13959_));
 NOR2_X2 _23656_ (.A1(_11062_),
    .A2(_17085_),
    .ZN(_13960_));
 CLKBUF_X2 _23657_ (.A(_13960_),
    .Z(_13961_));
 BUF_X2 _23658_ (.A(_13961_),
    .Z(_13962_));
 OAI21_X1 _23659_ (.A(_13953_),
    .B1(_13959_),
    .B2(_13962_),
    .ZN(_13963_));
 INV_X1 _23660_ (.A(_17088_),
    .ZN(_13964_));
 AND2_X1 _23661_ (.A1(_13964_),
    .A2(_17087_),
    .ZN(_13965_));
 AND2_X1 _23662_ (.A1(_13965_),
    .A2(_13950_),
    .ZN(_13966_));
 CLKBUF_X2 _23663_ (.A(_13966_),
    .Z(_13967_));
 INV_X1 _23664_ (.A(_13967_),
    .ZN(_13968_));
 INV_X1 _23665_ (.A(_17085_),
    .ZN(_13969_));
 NOR2_X2 _23666_ (.A1(_13969_),
    .A2(_17086_),
    .ZN(_13970_));
 INV_X1 _23667_ (.A(_17083_),
    .ZN(_13971_));
 NOR2_X1 _23668_ (.A1(_13971_),
    .A2(_11046_),
    .ZN(_13972_));
 BUF_X2 _23669_ (.A(_13972_),
    .Z(_13973_));
 AND2_X1 _23670_ (.A1(_13970_),
    .A2(_13973_),
    .ZN(_13974_));
 INV_X1 _23671_ (.A(_13974_),
    .ZN(_13975_));
 NOR2_X1 _23672_ (.A1(_17085_),
    .A2(_17086_),
    .ZN(_13976_));
 CLKBUF_X2 _23673_ (.A(_13976_),
    .Z(_13977_));
 AND2_X2 _23674_ (.A1(_13955_),
    .A2(_13977_),
    .ZN(_13978_));
 INV_X1 _23675_ (.A(_13978_),
    .ZN(_13979_));
 AOI21_X1 _23676_ (.A(_13968_),
    .B1(_13975_),
    .B2(_13979_),
    .ZN(_13980_));
 AND2_X1 _23677_ (.A1(_13960_),
    .A2(_17083_),
    .ZN(_13981_));
 NOR2_X1 _23678_ (.A1(_17087_),
    .A2(_17088_),
    .ZN(_13982_));
 CLKBUF_X2 _23679_ (.A(_13982_),
    .Z(_13983_));
 AND2_X1 _23680_ (.A1(_13950_),
    .A2(_13983_),
    .ZN(_13984_));
 NAND2_X1 _23681_ (.A1(_13981_),
    .A2(_13984_),
    .ZN(_13985_));
 NAND4_X1 _23682_ (.A1(_13955_),
    .A2(_13957_),
    .A3(_13950_),
    .A4(_13983_),
    .ZN(_13986_));
 AND2_X1 _23683_ (.A1(_13956_),
    .A2(_13954_),
    .ZN(_13987_));
 BUF_X2 _23684_ (.A(_13987_),
    .Z(_13988_));
 INV_X1 _23685_ (.A(_13988_),
    .ZN(_13989_));
 INV_X1 _23686_ (.A(_13984_),
    .ZN(_13990_));
 OAI211_X1 _23687_ (.A(_13985_),
    .B(_13986_),
    .C1(_13989_),
    .C2(_13990_),
    .ZN(_13991_));
 AND3_X1 _23688_ (.A1(_13984_),
    .A2(_13955_),
    .A3(_13977_),
    .ZN(_13992_));
 OR2_X1 _23689_ (.A1(_13991_),
    .A2(_13992_),
    .ZN(_13993_));
 BUF_X2 _23690_ (.A(_13966_),
    .Z(_13994_));
 INV_X1 _23691_ (.A(_13961_),
    .ZN(_13995_));
 NOR2_X2 _23692_ (.A1(_17083_),
    .A2(_17084_),
    .ZN(_13996_));
 INV_X1 _23693_ (.A(_13996_),
    .ZN(_13997_));
 NAND2_X1 _23694_ (.A1(_13997_),
    .A2(_13957_),
    .ZN(_13998_));
 AND2_X1 _23695_ (.A1(_17083_),
    .A2(_17084_),
    .ZN(_13999_));
 CLKBUF_X2 _23696_ (.A(_13999_),
    .Z(_14000_));
 OAI21_X1 _23697_ (.A(_13995_),
    .B1(_13998_),
    .B2(_14000_),
    .ZN(_14001_));
 AOI211_X1 _23698_ (.A(_13980_),
    .B(_13993_),
    .C1(_13994_),
    .C2(_14001_),
    .ZN(_14002_));
 INV_X1 _23699_ (.A(_13955_),
    .ZN(_14003_));
 NOR2_X2 _23700_ (.A1(_13964_),
    .A2(_17087_),
    .ZN(_14004_));
 AND2_X1 _23701_ (.A1(_14004_),
    .A2(_13950_),
    .ZN(_14005_));
 BUF_X1 _23702_ (.A(_14005_),
    .Z(_14006_));
 INV_X1 _23703_ (.A(_13972_),
    .ZN(_14007_));
 BUF_X2 _23704_ (.A(_13977_),
    .Z(_14008_));
 AND4_X1 _23705_ (.A1(_14003_),
    .A2(_14006_),
    .A3(_14007_),
    .A4(_14008_),
    .ZN(_14009_));
 INV_X1 _23706_ (.A(_14006_),
    .ZN(_14010_));
 NAND2_X1 _23707_ (.A1(_14007_),
    .A2(_13960_),
    .ZN(_14011_));
 NOR2_X1 _23708_ (.A1(_14010_),
    .A2(_14011_),
    .ZN(_14012_));
 AND2_X2 _23709_ (.A1(_13970_),
    .A2(_13954_),
    .ZN(_14013_));
 AND2_X1 _23710_ (.A1(_14013_),
    .A2(_14006_),
    .ZN(_14014_));
 AND2_X1 _23711_ (.A1(_13957_),
    .A2(_17083_),
    .ZN(_14015_));
 AND2_X1 _23712_ (.A1(_14006_),
    .A2(_14015_),
    .ZN(_14016_));
 NOR4_X1 _23713_ (.A1(_14009_),
    .A2(_14012_),
    .A3(_14014_),
    .A4(_14016_),
    .ZN(_14017_));
 AND2_X1 _23714_ (.A1(_13970_),
    .A2(_13996_),
    .ZN(_14018_));
 AND2_X1 _23715_ (.A1(_14018_),
    .A2(_13951_),
    .ZN(_14019_));
 AND2_X2 _23716_ (.A1(_13973_),
    .A2(_13977_),
    .ZN(_14020_));
 AND2_X1 _23717_ (.A1(_14020_),
    .A2(_13951_),
    .ZN(_14021_));
 AND2_X2 _23718_ (.A1(_13977_),
    .A2(_11046_),
    .ZN(_14022_));
 AOI211_X1 _23719_ (.A(_14019_),
    .B(_14021_),
    .C1(_14022_),
    .C2(_13953_),
    .ZN(_14023_));
 AND4_X1 _23720_ (.A1(_13963_),
    .A2(_14002_),
    .A3(_14017_),
    .A4(_14023_),
    .ZN(_14024_));
 AND2_X1 _23721_ (.A1(_13960_),
    .A2(_13996_),
    .ZN(_14025_));
 NOR2_X2 _23722_ (.A1(_17090_),
    .A2(_17091_),
    .ZN(_14026_));
 AND2_X1 _23723_ (.A1(_13949_),
    .A2(_14026_),
    .ZN(_14027_));
 AND2_X1 _23724_ (.A1(_14025_),
    .A2(_14027_),
    .ZN(_14028_));
 INV_X1 _23725_ (.A(_14027_),
    .ZN(_14029_));
 AND2_X1 _23726_ (.A1(_13956_),
    .A2(_13999_),
    .ZN(_14030_));
 BUF_X2 _23727_ (.A(_14030_),
    .Z(_14031_));
 INV_X1 _23728_ (.A(_14031_),
    .ZN(_14032_));
 AOI21_X1 _23729_ (.A(_14029_),
    .B1(_13989_),
    .B2(_14032_),
    .ZN(_14033_));
 NAND2_X1 _23730_ (.A1(_13997_),
    .A2(_13977_),
    .ZN(_14034_));
 NOR2_X1 _23731_ (.A1(_14029_),
    .A2(_14034_),
    .ZN(_14035_));
 CLKBUF_X2 _23732_ (.A(_13970_),
    .Z(_14036_));
 CLKBUF_X2 _23733_ (.A(_13955_),
    .Z(_14037_));
 AND3_X1 _23734_ (.A1(_14027_),
    .A2(_14036_),
    .A3(_14037_),
    .ZN(_14038_));
 OR4_X1 _23735_ (.A1(_14028_),
    .A2(_14033_),
    .A3(_14035_),
    .A4(_14038_),
    .ZN(_14039_));
 AND2_X1 _23736_ (.A1(_14026_),
    .A2(_13982_),
    .ZN(_14040_));
 BUF_X1 _23737_ (.A(_14040_),
    .Z(_14041_));
 AND2_X1 _23738_ (.A1(_13974_),
    .A2(_14041_),
    .ZN(_14042_));
 AND2_X2 _23739_ (.A1(_13970_),
    .A2(_11046_),
    .ZN(_14043_));
 AND2_X1 _23740_ (.A1(_14043_),
    .A2(_14041_),
    .ZN(_14044_));
 AND2_X1 _23741_ (.A1(_14041_),
    .A2(_14022_),
    .ZN(_14045_));
 NOR3_X1 _23742_ (.A1(_14042_),
    .A2(_14044_),
    .A3(_14045_),
    .ZN(_14046_));
 BUF_X2 _23743_ (.A(_14040_),
    .Z(_14047_));
 NAND3_X1 _23744_ (.A1(_14047_),
    .A2(_13997_),
    .A3(_13962_),
    .ZN(_14048_));
 INV_X1 _23745_ (.A(_14047_),
    .ZN(_14049_));
 NOR2_X1 _23746_ (.A1(_13998_),
    .A2(_14000_),
    .ZN(_14050_));
 INV_X1 _23747_ (.A(_14050_),
    .ZN(_14051_));
 OAI211_X1 _23748_ (.A(_14046_),
    .B(_14048_),
    .C1(_14049_),
    .C2(_14051_),
    .ZN(_14052_));
 AND2_X1 _23749_ (.A1(_13965_),
    .A2(_14026_),
    .ZN(_14053_));
 CLKBUF_X2 _23750_ (.A(_14053_),
    .Z(_14054_));
 AND2_X1 _23751_ (.A1(_14000_),
    .A2(_13977_),
    .ZN(_14055_));
 BUF_X2 _23752_ (.A(_14055_),
    .Z(_14056_));
 OAI21_X1 _23753_ (.A(_14054_),
    .B1(_13978_),
    .B2(_14056_),
    .ZN(_14057_));
 AND2_X1 _23754_ (.A1(_13960_),
    .A2(_14000_),
    .ZN(_14058_));
 BUF_X2 _23755_ (.A(_14058_),
    .Z(_14059_));
 OAI21_X1 _23756_ (.A(_14054_),
    .B1(_14025_),
    .B2(_14059_),
    .ZN(_14060_));
 INV_X2 _23757_ (.A(_13999_),
    .ZN(_14061_));
 NAND2_X1 _23758_ (.A1(_14061_),
    .A2(_14036_),
    .ZN(_14062_));
 NOR2_X1 _23759_ (.A1(_14062_),
    .A2(_13996_),
    .ZN(_14063_));
 INV_X1 _23760_ (.A(_14063_),
    .ZN(_14064_));
 INV_X1 _23761_ (.A(_14053_),
    .ZN(_14065_));
 OAI211_X1 _23762_ (.A(_14057_),
    .B(_14060_),
    .C1(_14064_),
    .C2(_14065_),
    .ZN(_14066_));
 AND2_X1 _23763_ (.A1(_14004_),
    .A2(_14026_),
    .ZN(_14067_));
 INV_X1 _23764_ (.A(_13977_),
    .ZN(_14068_));
 NOR2_X1 _23765_ (.A1(_14068_),
    .A2(_14000_),
    .ZN(_14069_));
 AND2_X1 _23766_ (.A1(_14067_),
    .A2(_14069_),
    .ZN(_14070_));
 INV_X1 _23767_ (.A(_14070_),
    .ZN(_14071_));
 NAND4_X1 _23768_ (.A1(_14067_),
    .A2(_13997_),
    .A3(_14061_),
    .A4(_14036_),
    .ZN(_14072_));
 AND2_X1 _23769_ (.A1(_13997_),
    .A2(_13960_),
    .ZN(_14073_));
 NAND2_X1 _23770_ (.A1(_14073_),
    .A2(_14067_),
    .ZN(_14074_));
 AND2_X1 _23771_ (.A1(_13957_),
    .A2(_13996_),
    .ZN(_14075_));
 CLKBUF_X2 _23772_ (.A(_14075_),
    .Z(_14076_));
 AND2_X1 _23773_ (.A1(_11046_),
    .A2(_17086_),
    .ZN(_14077_));
 AND2_X1 _23774_ (.A1(_14077_),
    .A2(_17085_),
    .ZN(_14078_));
 BUF_X2 _23775_ (.A(_14078_),
    .Z(_14079_));
 OAI21_X1 _23776_ (.A(_14067_),
    .B1(_14076_),
    .B2(_14079_),
    .ZN(_14080_));
 NAND4_X1 _23777_ (.A1(_14071_),
    .A2(_14072_),
    .A3(_14074_),
    .A4(_14080_),
    .ZN(_14081_));
 NOR4_X1 _23778_ (.A1(_14039_),
    .A2(_14052_),
    .A3(_14066_),
    .A4(_14081_),
    .ZN(_14082_));
 INV_X1 _23779_ (.A(_13998_),
    .ZN(_14083_));
 INV_X1 _23780_ (.A(_17090_),
    .ZN(_14084_));
 NOR2_X1 _23781_ (.A1(_14084_),
    .A2(_17091_),
    .ZN(_14085_));
 CLKBUF_X2 _23782_ (.A(_14085_),
    .Z(_14086_));
 AND2_X2 _23783_ (.A1(_14086_),
    .A2(_13949_),
    .ZN(_14087_));
 NAND3_X1 _23784_ (.A1(_14083_),
    .A2(_14061_),
    .A3(_14087_),
    .ZN(_14088_));
 NAND2_X1 _23785_ (.A1(_14059_),
    .A2(_14087_),
    .ZN(_14089_));
 AND2_X1 _23786_ (.A1(_14088_),
    .A2(_14089_),
    .ZN(_14090_));
 AND2_X2 _23787_ (.A1(_14004_),
    .A2(_14085_),
    .ZN(_14091_));
 AND2_X2 _23788_ (.A1(_13970_),
    .A2(_14000_),
    .ZN(_14092_));
 AND2_X1 _23789_ (.A1(_14091_),
    .A2(_14092_),
    .ZN(_14093_));
 INV_X1 _23790_ (.A(_14093_),
    .ZN(_14094_));
 AND2_X1 _23791_ (.A1(_13970_),
    .A2(_13955_),
    .ZN(_14095_));
 NAND2_X1 _23792_ (.A1(_14095_),
    .A2(_14091_),
    .ZN(_14096_));
 INV_X1 _23793_ (.A(_14013_),
    .ZN(_14097_));
 INV_X1 _23794_ (.A(_14091_),
    .ZN(_14098_));
 OAI211_X1 _23795_ (.A(_14094_),
    .B(_14096_),
    .C1(_14097_),
    .C2(_14098_),
    .ZN(_14099_));
 BUF_X2 _23796_ (.A(_13954_),
    .Z(_14100_));
 OAI21_X1 _23797_ (.A(_13961_),
    .B1(_17083_),
    .B2(_14100_),
    .ZN(_14101_));
 NOR2_X1 _23798_ (.A1(_14098_),
    .A2(_14101_),
    .ZN(_14102_));
 NAND2_X1 _23799_ (.A1(_14091_),
    .A2(_14020_),
    .ZN(_14103_));
 INV_X1 _23800_ (.A(_14055_),
    .ZN(_14104_));
 OAI21_X1 _23801_ (.A(_14103_),
    .B1(_14098_),
    .B2(_14104_),
    .ZN(_14105_));
 AND2_X1 _23802_ (.A1(_14091_),
    .A2(_13959_),
    .ZN(_14106_));
 NOR4_X1 _23803_ (.A1(_14099_),
    .A2(_14102_),
    .A3(_14105_),
    .A4(_14106_),
    .ZN(_14107_));
 AND2_X1 _23804_ (.A1(_13965_),
    .A2(_14086_),
    .ZN(_14108_));
 INV_X1 _23805_ (.A(_14108_),
    .ZN(_14109_));
 INV_X1 _23806_ (.A(_13981_),
    .ZN(_14110_));
 AOI21_X1 _23807_ (.A(_14109_),
    .B1(_14032_),
    .B2(_14110_),
    .ZN(_14111_));
 INV_X1 _23808_ (.A(_14043_),
    .ZN(_14112_));
 NAND2_X2 _23809_ (.A1(_14003_),
    .A2(_14008_),
    .ZN(_14113_));
 AOI21_X1 _23810_ (.A(_14109_),
    .B1(_14112_),
    .B2(_14113_),
    .ZN(_14114_));
 AND2_X1 _23811_ (.A1(_14086_),
    .A2(_13983_),
    .ZN(_14115_));
 INV_X1 _23812_ (.A(_14115_),
    .ZN(_14116_));
 INV_X1 _23813_ (.A(_14018_),
    .ZN(_14117_));
 AND2_X2 _23814_ (.A1(_13977_),
    .A2(_13954_),
    .ZN(_14118_));
 INV_X2 _23815_ (.A(_14118_),
    .ZN(_14119_));
 AOI21_X1 _23816_ (.A(_14116_),
    .B1(_14117_),
    .B2(_14119_),
    .ZN(_14120_));
 OAI21_X1 _23817_ (.A(_14115_),
    .B1(_13959_),
    .B2(_13988_),
    .ZN(_14121_));
 NAND4_X1 _23818_ (.A1(_13961_),
    .A2(_14086_),
    .A3(_11039_),
    .A4(_13983_),
    .ZN(_14122_));
 NAND2_X1 _23819_ (.A1(_14121_),
    .A2(_14122_),
    .ZN(_14123_));
 NOR4_X1 _23820_ (.A1(_14111_),
    .A2(_14114_),
    .A3(_14120_),
    .A4(_14123_),
    .ZN(_14124_));
 AND2_X1 _23821_ (.A1(_14087_),
    .A2(_14055_),
    .ZN(_14125_));
 NAND2_X1 _23822_ (.A1(_14020_),
    .A2(_14087_),
    .ZN(_14126_));
 INV_X1 _23823_ (.A(_14087_),
    .ZN(_14127_));
 AND2_X1 _23824_ (.A1(_13996_),
    .A2(_13976_),
    .ZN(_14128_));
 BUF_X2 _23825_ (.A(_14128_),
    .Z(_14129_));
 INV_X1 _23826_ (.A(_14129_),
    .ZN(_14130_));
 OAI21_X1 _23827_ (.A(_14126_),
    .B1(_14127_),
    .B2(_14130_),
    .ZN(_14131_));
 AND2_X2 _23828_ (.A1(_14036_),
    .A2(_11039_),
    .ZN(_14132_));
 BUF_X2 _23829_ (.A(_14087_),
    .Z(_14133_));
 AOI211_X1 _23830_ (.A(_14125_),
    .B(_14131_),
    .C1(_14132_),
    .C2(_14133_),
    .ZN(_14134_));
 AND4_X1 _23831_ (.A1(_14090_),
    .A2(_14107_),
    .A3(_14124_),
    .A4(_14134_),
    .ZN(_14135_));
 AND2_X1 _23832_ (.A1(_14084_),
    .A2(_17091_),
    .ZN(_14136_));
 AND2_X2 _23833_ (.A1(_13965_),
    .A2(_14136_),
    .ZN(_14137_));
 AND3_X1 _23834_ (.A1(_14137_),
    .A2(_13997_),
    .A3(_14069_),
    .ZN(_14138_));
 AOI21_X1 _23835_ (.A(_14138_),
    .B1(_14079_),
    .B2(_14137_),
    .ZN(_14139_));
 INV_X1 _23836_ (.A(_13970_),
    .ZN(_14140_));
 NOR2_X2 _23837_ (.A1(_14140_),
    .A2(_13955_),
    .ZN(_14141_));
 AND2_X1 _23838_ (.A1(_14136_),
    .A2(_13983_),
    .ZN(_14142_));
 BUF_X2 _23839_ (.A(_14142_),
    .Z(_14143_));
 NAND2_X1 _23840_ (.A1(_14141_),
    .A2(_14143_),
    .ZN(_14144_));
 BUF_X2 _23841_ (.A(_14136_),
    .Z(_14145_));
 BUF_X2 _23842_ (.A(_13971_),
    .Z(_14146_));
 NAND4_X1 _23843_ (.A1(_14145_),
    .A2(_14146_),
    .A3(_13983_),
    .A4(_14008_),
    .ZN(_14147_));
 OAI21_X1 _23844_ (.A(_14143_),
    .B1(_14083_),
    .B2(_13981_),
    .ZN(_14148_));
 NAND4_X1 _23845_ (.A1(_14139_),
    .A2(_14144_),
    .A3(_14147_),
    .A4(_14148_),
    .ZN(_14149_));
 OAI211_X1 _23846_ (.A(_14004_),
    .B(_14136_),
    .C1(_14031_),
    .C2(_13988_),
    .ZN(_14150_));
 NAND4_X1 _23847_ (.A1(_14145_),
    .A2(_14004_),
    .A3(_13961_),
    .A4(_13973_),
    .ZN(_14151_));
 NAND2_X1 _23848_ (.A1(_14150_),
    .A2(_14151_),
    .ZN(_14152_));
 AND2_X1 _23849_ (.A1(_14136_),
    .A2(_13949_),
    .ZN(_14153_));
 AND2_X1 _23850_ (.A1(_14141_),
    .A2(_14153_),
    .ZN(_14154_));
 NOR2_X1 _23851_ (.A1(_14068_),
    .A2(_13973_),
    .ZN(_14155_));
 AND2_X1 _23852_ (.A1(_14153_),
    .A2(_14155_),
    .ZN(_14156_));
 AND2_X1 _23853_ (.A1(_14153_),
    .A2(_14075_),
    .ZN(_14157_));
 OR3_X1 _23854_ (.A1(_14154_),
    .A2(_14156_),
    .A3(_14157_),
    .ZN(_14158_));
 AND2_X1 _23855_ (.A1(_14136_),
    .A2(_14004_),
    .ZN(_14159_));
 BUF_X2 _23856_ (.A(_14159_),
    .Z(_14160_));
 AND2_X1 _23857_ (.A1(_14160_),
    .A2(_14018_),
    .ZN(_14161_));
 NOR4_X1 _23858_ (.A1(_14149_),
    .A2(_14152_),
    .A3(_14158_),
    .A4(_14161_),
    .ZN(_14162_));
 NAND4_X1 _23859_ (.A1(_14024_),
    .A2(_14082_),
    .A3(_14135_),
    .A4(_14162_),
    .ZN(_14163_));
 AND2_X1 _23860_ (.A1(_14047_),
    .A2(_14129_),
    .ZN(_14164_));
 NOR2_X1 _23861_ (.A1(_14163_),
    .A2(_14164_),
    .ZN(_14165_));
 INV_X1 _23862_ (.A(_00988_),
    .ZN(_14166_));
 XNOR2_X1 _23863_ (.A(_14165_),
    .B(_14166_),
    .ZN(_14167_));
 MUX2_X1 _23864_ (.A(_01325_),
    .B(_14167_),
    .S(_03749_),
    .Z(_01058_));
 AND2_X1 _23865_ (.A1(_14153_),
    .A2(_13958_),
    .ZN(_14168_));
 AND2_X1 _23866_ (.A1(_14153_),
    .A2(_13987_),
    .ZN(_14169_));
 AOI221_X4 _23867_ (.A(_14168_),
    .B1(_14153_),
    .B2(_13981_),
    .C1(_11039_),
    .C2(_14169_),
    .ZN(_14170_));
 BUF_X2 _23868_ (.A(_14153_),
    .Z(_14171_));
 AND2_X1 _23869_ (.A1(_14008_),
    .A2(_14146_),
    .ZN(_14172_));
 OAI21_X1 _23870_ (.A(_14171_),
    .B1(_14095_),
    .B2(_14172_),
    .ZN(_14173_));
 AND2_X1 _23871_ (.A1(_14170_),
    .A2(_14173_),
    .ZN(_14174_));
 AND2_X1 _23872_ (.A1(_14159_),
    .A2(_14022_),
    .ZN(_14175_));
 AND2_X1 _23873_ (.A1(_14159_),
    .A2(_14020_),
    .ZN(_14176_));
 BUF_X2 _23874_ (.A(_13974_),
    .Z(_14177_));
 AOI211_X1 _23875_ (.A(_14175_),
    .B(_14176_),
    .C1(_14177_),
    .C2(_14160_),
    .ZN(_14178_));
 INV_X1 _23876_ (.A(_14159_),
    .ZN(_14179_));
 OAI211_X1 _23877_ (.A(_14174_),
    .B(_14178_),
    .C1(_14179_),
    .C2(_14101_),
    .ZN(_14180_));
 NAND4_X1 _23878_ (.A1(_14136_),
    .A2(_13983_),
    .A3(_14037_),
    .A4(_14008_),
    .ZN(_14181_));
 NAND2_X1 _23879_ (.A1(_14144_),
    .A2(_14181_),
    .ZN(_14182_));
 INV_X1 _23880_ (.A(_14142_),
    .ZN(_14183_));
 AND2_X1 _23881_ (.A1(_14073_),
    .A2(_14061_),
    .ZN(_14184_));
 INV_X1 _23882_ (.A(_14184_),
    .ZN(_14185_));
 AOI21_X1 _23883_ (.A(_14183_),
    .B1(_14185_),
    .B2(_14032_),
    .ZN(_14186_));
 INV_X1 _23884_ (.A(_14137_),
    .ZN(_14187_));
 AOI21_X1 _23885_ (.A(_14187_),
    .B1(_14097_),
    .B2(_13979_),
    .ZN(_14188_));
 AND2_X2 _23886_ (.A1(_13960_),
    .A2(_13954_),
    .ZN(_14189_));
 NAND2_X1 _23887_ (.A1(_14137_),
    .A2(_14189_),
    .ZN(_14190_));
 INV_X1 _23888_ (.A(_13957_),
    .ZN(_14191_));
 OAI21_X1 _23889_ (.A(_14190_),
    .B1(_14187_),
    .B2(_14191_),
    .ZN(_14192_));
 OR4_X1 _23890_ (.A1(_14182_),
    .A2(_14186_),
    .A3(_14188_),
    .A4(_14192_),
    .ZN(_14193_));
 CLKBUF_X2 _23891_ (.A(_13965_),
    .Z(_14194_));
 AND4_X1 _23892_ (.A1(_11039_),
    .A2(_14194_),
    .A3(_13950_),
    .A4(_13977_),
    .ZN(_14195_));
 AND2_X1 _23893_ (.A1(_13967_),
    .A2(_13974_),
    .ZN(_14196_));
 AOI211_X1 _23894_ (.A(_14195_),
    .B(_14196_),
    .C1(_14043_),
    .C2(_13994_),
    .ZN(_14197_));
 CLKBUF_X2 _23895_ (.A(_13984_),
    .Z(_14198_));
 BUF_X2 _23896_ (.A(_14198_),
    .Z(_14199_));
 NAND2_X1 _23897_ (.A1(_14104_),
    .A2(_14130_),
    .ZN(_14200_));
 OAI21_X1 _23898_ (.A(_14199_),
    .B1(_14200_),
    .B2(_14132_),
    .ZN(_14201_));
 AND2_X1 _23899_ (.A1(_14058_),
    .A2(_14198_),
    .ZN(_14202_));
 AND2_X1 _23900_ (.A1(_14078_),
    .A2(_14198_),
    .ZN(_14203_));
 AND2_X1 _23901_ (.A1(_14075_),
    .A2(_13984_),
    .ZN(_14204_));
 NOR3_X1 _23902_ (.A1(_14202_),
    .A2(_14203_),
    .A3(_14204_),
    .ZN(_14205_));
 AND2_X1 _23903_ (.A1(_13960_),
    .A2(_13955_),
    .ZN(_14206_));
 AND2_X1 _23904_ (.A1(_13967_),
    .A2(_14206_),
    .ZN(_14207_));
 INV_X1 _23905_ (.A(_14207_),
    .ZN(_14208_));
 OAI21_X1 _23906_ (.A(_13967_),
    .B1(_14076_),
    .B2(_14031_),
    .ZN(_14209_));
 AND2_X1 _23907_ (.A1(_14208_),
    .A2(_14209_),
    .ZN(_14210_));
 NAND4_X1 _23908_ (.A1(_14197_),
    .A2(_14201_),
    .A3(_14205_),
    .A4(_14210_),
    .ZN(_14211_));
 AND2_X1 _23909_ (.A1(_14005_),
    .A2(_14075_),
    .ZN(_14212_));
 AND3_X1 _23910_ (.A1(_14031_),
    .A2(_14004_),
    .A3(_13950_),
    .ZN(_14213_));
 OR2_X1 _23911_ (.A1(_14212_),
    .A2(_14213_),
    .ZN(_14214_));
 BUF_X2 _23912_ (.A(_14206_),
    .Z(_14215_));
 AND2_X1 _23913_ (.A1(_14215_),
    .A2(_14006_),
    .ZN(_14216_));
 AND2_X1 _23914_ (.A1(_14189_),
    .A2(_14006_),
    .ZN(_14217_));
 AND2_X1 _23915_ (.A1(_14095_),
    .A2(_14006_),
    .ZN(_14218_));
 NOR4_X1 _23916_ (.A1(_14214_),
    .A2(_14216_),
    .A3(_14217_),
    .A4(_14218_),
    .ZN(_14219_));
 NAND2_X1 _23917_ (.A1(_14013_),
    .A2(_13952_),
    .ZN(_14220_));
 NAND2_X1 _23918_ (.A1(_14095_),
    .A2(_13953_),
    .ZN(_14221_));
 OAI21_X1 _23919_ (.A(_13953_),
    .B1(_14059_),
    .B2(_14079_),
    .ZN(_14222_));
 NAND4_X1 _23920_ (.A1(_14219_),
    .A2(_14220_),
    .A3(_14221_),
    .A4(_14222_),
    .ZN(_14223_));
 NOR4_X1 _23921_ (.A1(_14180_),
    .A2(_14193_),
    .A3(_14211_),
    .A4(_14223_),
    .ZN(_14224_));
 BUF_X2 _23922_ (.A(_14054_),
    .Z(_14225_));
 AND2_X1 _23923_ (.A1(_14036_),
    .A2(_13971_),
    .ZN(_14226_));
 OAI21_X1 _23924_ (.A(_14225_),
    .B1(_14226_),
    .B2(_14118_),
    .ZN(_14227_));
 AND3_X1 _23925_ (.A1(_14040_),
    .A2(_13996_),
    .A3(_14036_),
    .ZN(_14228_));
 AND3_X1 _23926_ (.A1(_14041_),
    .A2(_14036_),
    .A3(_14037_),
    .ZN(_14229_));
 NOR4_X1 _23927_ (.A1(_14042_),
    .A2(_14228_),
    .A3(_14229_),
    .A4(_14045_),
    .ZN(_14230_));
 NAND3_X1 _23928_ (.A1(_14047_),
    .A2(_13962_),
    .A3(_14037_),
    .ZN(_14231_));
 OAI21_X1 _23929_ (.A(_14047_),
    .B1(_13959_),
    .B2(_14031_),
    .ZN(_14232_));
 NAND3_X1 _23930_ (.A1(_14047_),
    .A2(_14000_),
    .A3(_13962_),
    .ZN(_14233_));
 NAND2_X1 _23931_ (.A1(_13988_),
    .A2(_14047_),
    .ZN(_14234_));
 AND4_X1 _23932_ (.A1(_14231_),
    .A2(_14232_),
    .A3(_14233_),
    .A4(_14234_),
    .ZN(_14235_));
 AND2_X1 _23933_ (.A1(_14077_),
    .A2(_13969_),
    .ZN(_14236_));
 BUF_X2 _23934_ (.A(_14236_),
    .Z(_14237_));
 OAI21_X1 _23935_ (.A(_14225_),
    .B1(_13959_),
    .B2(_14237_),
    .ZN(_14238_));
 AND4_X1 _23936_ (.A1(_14227_),
    .A2(_14230_),
    .A3(_14235_),
    .A4(_14238_),
    .ZN(_14239_));
 NOR3_X1 _23937_ (.A1(_17087_),
    .A2(_17090_),
    .A3(_17091_),
    .ZN(_14240_));
 NAND3_X1 _23938_ (.A1(_14061_),
    .A2(_14240_),
    .A3(_13970_),
    .ZN(_14241_));
 NOR2_X1 _23939_ (.A1(_14241_),
    .A2(_13964_),
    .ZN(_14242_));
 INV_X1 _23940_ (.A(_14242_),
    .ZN(_14243_));
 INV_X1 _23941_ (.A(_13959_),
    .ZN(_14244_));
 AOI21_X1 _23942_ (.A(_14029_),
    .B1(_14244_),
    .B2(_13989_),
    .ZN(_14245_));
 AND2_X1 _23943_ (.A1(_13960_),
    .A2(_13973_),
    .ZN(_14246_));
 AND2_X1 _23944_ (.A1(_14246_),
    .A2(_14027_),
    .ZN(_14247_));
 AND2_X1 _23945_ (.A1(_14058_),
    .A2(_14027_),
    .ZN(_14248_));
 NOR4_X1 _23946_ (.A1(_14245_),
    .A2(_14028_),
    .A3(_14247_),
    .A4(_14248_),
    .ZN(_14249_));
 BUF_X2 _23947_ (.A(_14067_),
    .Z(_14250_));
 NAND2_X1 _23948_ (.A1(_14250_),
    .A2(_14155_),
    .ZN(_14251_));
 CLKBUF_X2 _23949_ (.A(_14027_),
    .Z(_14252_));
 INV_X1 _23950_ (.A(_14034_),
    .ZN(_14253_));
 OAI21_X1 _23951_ (.A(_14252_),
    .B1(_14253_),
    .B2(_14132_),
    .ZN(_14254_));
 AND4_X1 _23952_ (.A1(_14243_),
    .A2(_14249_),
    .A3(_14251_),
    .A4(_14254_),
    .ZN(_14255_));
 AND2_X1 _23953_ (.A1(_14108_),
    .A2(_14189_),
    .ZN(_14256_));
 INV_X1 _23954_ (.A(_14256_),
    .ZN(_14257_));
 BUF_X2 _23955_ (.A(_14108_),
    .Z(_14258_));
 OAI21_X1 _23956_ (.A(_14258_),
    .B1(_14092_),
    .B2(_14129_),
    .ZN(_14259_));
 NAND3_X1 _23957_ (.A1(_14215_),
    .A2(_14194_),
    .A3(_14086_),
    .ZN(_14260_));
 OAI211_X1 _23958_ (.A(_14194_),
    .B(_14086_),
    .C1(_14031_),
    .C2(_14076_),
    .ZN(_14261_));
 NAND4_X1 _23959_ (.A1(_14257_),
    .A2(_14259_),
    .A3(_14260_),
    .A4(_14261_),
    .ZN(_14262_));
 BUF_X2 _23960_ (.A(_14115_),
    .Z(_14263_));
 INV_X1 _23961_ (.A(_14062_),
    .ZN(_14264_));
 AND2_X1 _23962_ (.A1(_14008_),
    .A2(_11039_),
    .ZN(_14265_));
 OAI21_X1 _23963_ (.A(_14263_),
    .B1(_14264_),
    .B2(_14265_),
    .ZN(_14266_));
 BUF_X2 _23964_ (.A(_13957_),
    .Z(_14267_));
 OAI211_X1 _23965_ (.A(_14263_),
    .B(_14267_),
    .C1(_14037_),
    .C2(_13973_),
    .ZN(_14268_));
 OAI211_X1 _23966_ (.A(_14266_),
    .B(_14268_),
    .C1(_13995_),
    .C2(_14116_),
    .ZN(_14269_));
 BUF_X2 _23967_ (.A(_14091_),
    .Z(_14270_));
 OAI21_X1 _23968_ (.A(_14270_),
    .B1(_13959_),
    .B2(_14237_),
    .ZN(_14271_));
 NAND2_X1 _23969_ (.A1(_14253_),
    .A2(_14270_),
    .ZN(_14272_));
 INV_X1 _23970_ (.A(_14226_),
    .ZN(_14273_));
 OAI211_X1 _23971_ (.A(_14271_),
    .B(_14272_),
    .C1(_14273_),
    .C2(_14098_),
    .ZN(_14274_));
 OAI21_X1 _23972_ (.A(_14087_),
    .B1(_14020_),
    .B2(_14056_),
    .ZN(_14275_));
 NAND3_X1 _23973_ (.A1(_14073_),
    .A2(_14133_),
    .A3(_14061_),
    .ZN(_14276_));
 NAND2_X1 _23974_ (.A1(_14083_),
    .A2(_14133_),
    .ZN(_14277_));
 CLKBUF_X2 _23975_ (.A(_14036_),
    .Z(_14278_));
 NAND4_X1 _23976_ (.A1(_14278_),
    .A2(_14086_),
    .A3(_13996_),
    .A4(_13949_),
    .ZN(_14279_));
 NAND4_X1 _23977_ (.A1(_14275_),
    .A2(_14276_),
    .A3(_14277_),
    .A4(_14279_),
    .ZN(_14280_));
 NOR4_X1 _23978_ (.A1(_14262_),
    .A2(_14269_),
    .A3(_14274_),
    .A4(_14280_),
    .ZN(_14281_));
 NAND4_X1 _23979_ (.A1(_14224_),
    .A2(_14239_),
    .A3(_14255_),
    .A4(_14281_),
    .ZN(_14282_));
 NOR2_X1 _23980_ (.A1(_14282_),
    .A2(_14164_),
    .ZN(_14283_));
 XOR2_X1 _23981_ (.A(_14283_),
    .B(_00989_),
    .Z(_14284_));
 BUF_X2 _23982_ (.A(_03738_),
    .Z(_14285_));
 MUX2_X1 _23983_ (.A(_01326_),
    .B(_14284_),
    .S(_14285_),
    .Z(_01069_));
 XOR2_X1 _23984_ (.A(_17193_),
    .B(_16997_),
    .Z(_14286_));
 XNOR2_X1 _23985_ (.A(_11312_),
    .B(_11776_),
    .ZN(_14287_));
 XOR2_X1 _23986_ (.A(_13842_),
    .B(_00990_),
    .Z(_14288_));
 XNOR2_X1 _23987_ (.A(_14287_),
    .B(_14288_),
    .ZN(_14289_));
 XOR2_X1 _23988_ (.A(_14289_),
    .B(_12500_),
    .Z(_14290_));
 MUX2_X1 _23989_ (.A(_14286_),
    .B(_14290_),
    .S(_11084_),
    .Z(_00684_));
 OAI21_X1 _23990_ (.A(_14198_),
    .B1(_14215_),
    .B2(_13981_),
    .ZN(_14291_));
 NAND3_X1 _23991_ (.A1(_13988_),
    .A2(_14198_),
    .A3(_11039_),
    .ZN(_14292_));
 AND2_X1 _23992_ (.A1(_14291_),
    .A2(_14292_),
    .ZN(_14293_));
 AND2_X1 _23993_ (.A1(_13966_),
    .A2(_14078_),
    .ZN(_14294_));
 AND2_X1 _23994_ (.A1(_13994_),
    .A2(_14076_),
    .ZN(_14295_));
 AND2_X1 _23995_ (.A1(_13967_),
    .A2(_14246_),
    .ZN(_14296_));
 NOR4_X1 _23996_ (.A1(_14207_),
    .A2(_14294_),
    .A3(_14295_),
    .A4(_14296_),
    .ZN(_14297_));
 AND2_X1 _23997_ (.A1(_14198_),
    .A2(_14055_),
    .ZN(_14298_));
 AOI211_X1 _23998_ (.A(_14298_),
    .B(_13992_),
    .C1(_14278_),
    .C2(_14199_),
    .ZN(_14299_));
 AND3_X1 _23999_ (.A1(_14020_),
    .A2(_14194_),
    .A3(_13950_),
    .ZN(_14300_));
 AND2_X1 _24000_ (.A1(_13967_),
    .A2(_14043_),
    .ZN(_14301_));
 AOI211_X1 _24001_ (.A(_14300_),
    .B(_14301_),
    .C1(_14022_),
    .C2(_13994_),
    .ZN(_14302_));
 AND4_X1 _24002_ (.A1(_14293_),
    .A2(_14297_),
    .A3(_14299_),
    .A4(_14302_),
    .ZN(_14303_));
 AOI21_X1 _24003_ (.A(_14183_),
    .B1(_13989_),
    .B2(_13995_),
    .ZN(_14304_));
 NAND3_X1 _24004_ (.A1(_14059_),
    .A2(_14194_),
    .A3(_14145_),
    .ZN(_14305_));
 OAI211_X1 _24005_ (.A(_14190_),
    .B(_14305_),
    .C1(_14187_),
    .C2(_13989_),
    .ZN(_14306_));
 AOI21_X1 _24006_ (.A(_14183_),
    .B1(_14140_),
    .B2(_14113_),
    .ZN(_14307_));
 AND2_X1 _24007_ (.A1(_14137_),
    .A2(_14022_),
    .ZN(_14308_));
 NOR4_X1 _24008_ (.A1(_14304_),
    .A2(_14306_),
    .A3(_14307_),
    .A4(_14308_),
    .ZN(_14309_));
 AND2_X1 _24009_ (.A1(_14043_),
    .A2(_14006_),
    .ZN(_14310_));
 INV_X1 _24010_ (.A(_14310_),
    .ZN(_14311_));
 INV_X1 _24011_ (.A(_13952_),
    .ZN(_14312_));
 INV_X1 _24012_ (.A(_14215_),
    .ZN(_14313_));
 INV_X1 _24013_ (.A(_14059_),
    .ZN(_14314_));
 AOI21_X1 _24014_ (.A(_14312_),
    .B1(_14313_),
    .B2(_14314_),
    .ZN(_14315_));
 AOI21_X1 _24015_ (.A(_14315_),
    .B1(_14015_),
    .B2(_13953_),
    .ZN(_14316_));
 BUF_X2 _24016_ (.A(_14005_),
    .Z(_14317_));
 NAND2_X1 _24017_ (.A1(_14003_),
    .A2(_13957_),
    .ZN(_14318_));
 INV_X1 _24018_ (.A(_14318_),
    .ZN(_14319_));
 OAI21_X1 _24019_ (.A(_14317_),
    .B1(_14184_),
    .B2(_14319_),
    .ZN(_14320_));
 OAI21_X1 _24020_ (.A(_13953_),
    .B1(_14200_),
    .B2(_14013_),
    .ZN(_14321_));
 AND4_X1 _24021_ (.A1(_14311_),
    .A2(_14316_),
    .A3(_14320_),
    .A4(_14321_),
    .ZN(_14322_));
 OAI21_X1 _24022_ (.A(_14160_),
    .B1(_14177_),
    .B2(_14043_),
    .ZN(_14323_));
 INV_X1 _24023_ (.A(_14153_),
    .ZN(_14324_));
 INV_X1 _24024_ (.A(_14189_),
    .ZN(_14325_));
 AOI21_X1 _24025_ (.A(_14324_),
    .B1(_14313_),
    .B2(_14325_),
    .ZN(_14326_));
 NOR3_X1 _24026_ (.A1(_14326_),
    .A2(_14157_),
    .A3(_14168_),
    .ZN(_14327_));
 OAI21_X1 _24027_ (.A(_14160_),
    .B1(_14050_),
    .B2(_14215_),
    .ZN(_14328_));
 OAI21_X1 _24028_ (.A(_14171_),
    .B1(_14264_),
    .B2(_14155_),
    .ZN(_14329_));
 AND4_X1 _24029_ (.A1(_14323_),
    .A2(_14327_),
    .A3(_14328_),
    .A4(_14329_),
    .ZN(_14330_));
 NAND4_X1 _24030_ (.A1(_14303_),
    .A2(_14309_),
    .A3(_14322_),
    .A4(_14330_),
    .ZN(_14331_));
 NOR2_X1 _24031_ (.A1(_14011_),
    .A2(_14037_),
    .ZN(_14332_));
 OAI21_X1 _24032_ (.A(_14270_),
    .B1(_14332_),
    .B2(_14050_),
    .ZN(_14333_));
 NAND2_X1 _24033_ (.A1(_14177_),
    .A2(_14270_),
    .ZN(_14334_));
 AND3_X1 _24034_ (.A1(_14094_),
    .A2(_14103_),
    .A3(_14334_),
    .ZN(_14335_));
 OAI21_X1 _24035_ (.A(_14133_),
    .B1(_14132_),
    .B2(_14056_),
    .ZN(_14336_));
 OAI211_X1 _24036_ (.A(_14133_),
    .B(_14100_),
    .C1(_14015_),
    .C2(_13962_),
    .ZN(_14337_));
 AND4_X1 _24037_ (.A1(_14333_),
    .A2(_14335_),
    .A3(_14336_),
    .A4(_14337_),
    .ZN(_14338_));
 AND3_X1 _24038_ (.A1(_14041_),
    .A2(_13961_),
    .A3(_14037_),
    .ZN(_14339_));
 AND3_X1 _24039_ (.A1(_14041_),
    .A2(_13957_),
    .A3(_14003_),
    .ZN(_14340_));
 OR2_X1 _24040_ (.A1(_14339_),
    .A2(_14340_),
    .ZN(_14341_));
 NAND2_X1 _24041_ (.A1(_14253_),
    .A2(_14041_),
    .ZN(_14342_));
 OAI22_X1 _24042_ (.A1(_14342_),
    .A2(_14000_),
    .B1(_14049_),
    .B2(_14112_),
    .ZN(_14343_));
 NAND2_X1 _24043_ (.A1(_14225_),
    .A2(_14059_),
    .ZN(_14344_));
 NAND2_X1 _24044_ (.A1(_14225_),
    .A2(_14189_),
    .ZN(_14345_));
 NAND2_X1 _24045_ (.A1(_14225_),
    .A2(_13988_),
    .ZN(_14346_));
 NAND3_X1 _24046_ (.A1(_14344_),
    .A2(_14345_),
    .A3(_14346_),
    .ZN(_14347_));
 NAND2_X1 _24047_ (.A1(_14054_),
    .A2(_14095_),
    .ZN(_14348_));
 OAI21_X1 _24048_ (.A(_14348_),
    .B1(_14065_),
    .B2(_14104_),
    .ZN(_14349_));
 NOR4_X1 _24049_ (.A1(_14341_),
    .A2(_14343_),
    .A3(_14347_),
    .A4(_14349_),
    .ZN(_14350_));
 AOI21_X1 _24050_ (.A(_14029_),
    .B1(_14064_),
    .B2(_14119_),
    .ZN(_14351_));
 AND4_X1 _24051_ (.A1(_11039_),
    .A2(_14267_),
    .A3(_13949_),
    .A4(_14026_),
    .ZN(_14352_));
 OR2_X1 _24052_ (.A1(_14028_),
    .A2(_14352_),
    .ZN(_14353_));
 NAND2_X1 _24053_ (.A1(_14250_),
    .A2(_14013_),
    .ZN(_14354_));
 NAND2_X1 _24054_ (.A1(_14250_),
    .A2(_14043_),
    .ZN(_14355_));
 INV_X1 _24055_ (.A(_14250_),
    .ZN(_14356_));
 OAI211_X1 _24056_ (.A(_14354_),
    .B(_14355_),
    .C1(_14356_),
    .C2(_14113_),
    .ZN(_14357_));
 NAND4_X1 _24057_ (.A1(_14004_),
    .A2(_13962_),
    .A3(_14037_),
    .A4(_14026_),
    .ZN(_14358_));
 NAND4_X1 _24058_ (.A1(_14004_),
    .A2(_14267_),
    .A3(_14000_),
    .A4(_14026_),
    .ZN(_14359_));
 OAI211_X1 _24059_ (.A(_14358_),
    .B(_14359_),
    .C1(_14356_),
    .C2(_14325_),
    .ZN(_14360_));
 NOR4_X1 _24060_ (.A1(_14351_),
    .A2(_14353_),
    .A3(_14357_),
    .A4(_14360_),
    .ZN(_14361_));
 OAI21_X1 _24061_ (.A(_14263_),
    .B1(_14177_),
    .B2(_13978_),
    .ZN(_14362_));
 OAI21_X1 _24062_ (.A(_14258_),
    .B1(_14177_),
    .B2(_14056_),
    .ZN(_14363_));
 OAI21_X1 _24063_ (.A(_14258_),
    .B1(_14215_),
    .B2(_14015_),
    .ZN(_14364_));
 OAI21_X1 _24064_ (.A(_14263_),
    .B1(_14215_),
    .B2(_14079_),
    .ZN(_14365_));
 AND4_X1 _24065_ (.A1(_14362_),
    .A2(_14363_),
    .A3(_14364_),
    .A4(_14365_),
    .ZN(_14366_));
 NAND4_X1 _24066_ (.A1(_14338_),
    .A2(_14350_),
    .A3(_14361_),
    .A4(_14366_),
    .ZN(_14367_));
 NOR2_X1 _24067_ (.A1(_14331_),
    .A2(_14367_),
    .ZN(_14368_));
 XOR2_X1 _24068_ (.A(_14368_),
    .B(_00991_),
    .Z(_14369_));
 MUX2_X1 _24069_ (.A(_01327_),
    .B(_14369_),
    .S(_14285_),
    .Z(_01080_));
 NAND4_X1 _24070_ (.A1(_14145_),
    .A2(_11040_),
    .A3(_13949_),
    .A4(_14008_),
    .ZN(_14370_));
 AND4_X1 _24071_ (.A1(_13961_),
    .A2(_14153_),
    .A3(_14003_),
    .A4(_14007_),
    .ZN(_14371_));
 AOI221_X4 _24072_ (.A(_14371_),
    .B1(_11039_),
    .B2(_14169_),
    .C1(_14079_),
    .C2(_14171_),
    .ZN(_14372_));
 OAI211_X1 _24073_ (.A(_14171_),
    .B(_14278_),
    .C1(_14146_),
    .C2(_11046_),
    .ZN(_14373_));
 AOI21_X1 _24074_ (.A(_14179_),
    .B1(_14032_),
    .B2(_14313_),
    .ZN(_14374_));
 AND2_X1 _24075_ (.A1(_14159_),
    .A2(_14092_),
    .ZN(_14375_));
 NOR4_X1 _24076_ (.A1(_14374_),
    .A2(_14161_),
    .A3(_14175_),
    .A4(_14375_),
    .ZN(_14376_));
 AND4_X1 _24077_ (.A1(_14370_),
    .A2(_14372_),
    .A3(_14373_),
    .A4(_14376_),
    .ZN(_14377_));
 AND2_X1 _24078_ (.A1(_14143_),
    .A2(_14237_),
    .ZN(_14378_));
 AOI21_X1 _24079_ (.A(_14183_),
    .B1(_14117_),
    .B2(_14113_),
    .ZN(_14379_));
 AOI211_X1 _24080_ (.A(_14378_),
    .B(_14379_),
    .C1(_14050_),
    .C2(_14143_),
    .ZN(_14380_));
 AOI21_X1 _24081_ (.A(_14187_),
    .B1(_14185_),
    .B2(_14191_),
    .ZN(_14381_));
 AOI211_X1 _24082_ (.A(_14308_),
    .B(_14381_),
    .C1(_14132_),
    .C2(_14137_),
    .ZN(_14382_));
 NAND2_X1 _24083_ (.A1(_14018_),
    .A2(_14199_),
    .ZN(_14383_));
 OAI21_X1 _24084_ (.A(_14198_),
    .B1(_13988_),
    .B2(_14078_),
    .ZN(_14384_));
 OAI211_X1 _24085_ (.A(_14198_),
    .B(_13962_),
    .C1(_11040_),
    .C2(_14100_),
    .ZN(_14385_));
 OAI21_X1 _24086_ (.A(_14198_),
    .B1(_14056_),
    .B2(_14118_),
    .ZN(_14386_));
 AND4_X1 _24087_ (.A1(_14383_),
    .A2(_14384_),
    .A3(_14385_),
    .A4(_14386_),
    .ZN(_14387_));
 AND3_X1 _24088_ (.A1(_14141_),
    .A2(_13994_),
    .A3(_14007_),
    .ZN(_14388_));
 AND2_X1 _24089_ (.A1(_13967_),
    .A2(_14058_),
    .ZN(_14389_));
 NOR4_X1 _24090_ (.A1(_14388_),
    .A2(_14389_),
    .A3(_14294_),
    .A4(_14300_),
    .ZN(_14390_));
 OAI211_X1 _24091_ (.A(_14317_),
    .B(_14008_),
    .C1(_14037_),
    .C2(_13973_),
    .ZN(_14391_));
 OAI211_X1 _24092_ (.A(_14317_),
    .B(_14036_),
    .C1(_14146_),
    .C2(_14100_),
    .ZN(_14392_));
 OAI211_X1 _24093_ (.A(_14317_),
    .B(_13961_),
    .C1(_11040_),
    .C2(_14100_),
    .ZN(_14393_));
 OAI21_X1 _24094_ (.A(_14317_),
    .B1(_14076_),
    .B2(_14078_),
    .ZN(_14394_));
 AND4_X1 _24095_ (.A1(_14391_),
    .A2(_14392_),
    .A3(_14393_),
    .A4(_14394_),
    .ZN(_14395_));
 NAND3_X1 _24096_ (.A1(_13952_),
    .A2(_14267_),
    .A3(_14037_),
    .ZN(_14396_));
 OAI211_X1 _24097_ (.A(_13952_),
    .B(_14036_),
    .C1(_13996_),
    .C2(_14000_),
    .ZN(_14397_));
 OAI211_X1 _24098_ (.A(_13952_),
    .B(_13961_),
    .C1(_11040_),
    .C2(_11046_),
    .ZN(_14398_));
 OAI21_X1 _24099_ (.A(_13952_),
    .B1(_14129_),
    .B2(_14022_),
    .ZN(_14399_));
 AND4_X1 _24100_ (.A1(_14396_),
    .A2(_14397_),
    .A3(_14398_),
    .A4(_14399_),
    .ZN(_14400_));
 AND4_X1 _24101_ (.A1(_14387_),
    .A2(_14390_),
    .A3(_14395_),
    .A4(_14400_),
    .ZN(_14401_));
 NAND4_X1 _24102_ (.A1(_14377_),
    .A2(_14380_),
    .A3(_14382_),
    .A4(_14401_),
    .ZN(_14402_));
 OAI21_X1 _24103_ (.A(_14047_),
    .B1(_14063_),
    .B2(_14265_),
    .ZN(_14403_));
 AND2_X1 _24104_ (.A1(_14076_),
    .A2(_14041_),
    .ZN(_14404_));
 AND2_X1 _24105_ (.A1(_13959_),
    .A2(_14041_),
    .ZN(_14405_));
 AOI211_X1 _24106_ (.A(_14404_),
    .B(_14405_),
    .C1(_14047_),
    .C2(_14059_),
    .ZN(_14406_));
 OAI21_X1 _24107_ (.A(_14225_),
    .B1(_14013_),
    .B2(_14155_),
    .ZN(_14407_));
 NAND2_X1 _24108_ (.A1(_14225_),
    .A2(_14076_),
    .ZN(_14408_));
 AND2_X1 _24109_ (.A1(_14060_),
    .A2(_14408_),
    .ZN(_14409_));
 AND4_X1 _24110_ (.A1(_14403_),
    .A2(_14406_),
    .A3(_14407_),
    .A4(_14409_),
    .ZN(_14410_));
 NAND2_X1 _24111_ (.A1(_14258_),
    .A2(_14267_),
    .ZN(_14411_));
 INV_X1 _24112_ (.A(_14237_),
    .ZN(_14412_));
 OAI211_X1 _24113_ (.A(_14257_),
    .B(_14411_),
    .C1(_14109_),
    .C2(_14412_),
    .ZN(_14413_));
 OAI211_X1 _24114_ (.A(_14263_),
    .B(_14008_),
    .C1(_14146_),
    .C2(_11046_),
    .ZN(_14414_));
 OAI21_X1 _24115_ (.A(_14414_),
    .B1(_14062_),
    .B2(_14116_),
    .ZN(_14415_));
 INV_X1 _24116_ (.A(_14246_),
    .ZN(_14416_));
 AND2_X1 _24117_ (.A1(_13957_),
    .A2(_13971_),
    .ZN(_14417_));
 INV_X1 _24118_ (.A(_14417_),
    .ZN(_14418_));
 AOI21_X1 _24119_ (.A(_14116_),
    .B1(_14416_),
    .B2(_14418_),
    .ZN(_14419_));
 INV_X1 _24120_ (.A(_14132_),
    .ZN(_14420_));
 AOI21_X1 _24121_ (.A(_14109_),
    .B1(_14420_),
    .B2(_14104_),
    .ZN(_14421_));
 NOR4_X1 _24122_ (.A1(_14413_),
    .A2(_14415_),
    .A3(_14419_),
    .A4(_14421_),
    .ZN(_14422_));
 AND2_X2 _24123_ (.A1(_13973_),
    .A2(_14267_),
    .ZN(_14423_));
 NAND2_X1 _24124_ (.A1(_14250_),
    .A2(_14423_),
    .ZN(_14424_));
 OAI21_X1 _24125_ (.A(_14250_),
    .B1(_14020_),
    .B2(_14132_),
    .ZN(_14425_));
 NAND3_X1 _24126_ (.A1(_14141_),
    .A2(_14252_),
    .A3(_14007_),
    .ZN(_14426_));
 NAND2_X1 _24127_ (.A1(_14076_),
    .A2(_14252_),
    .ZN(_14427_));
 AND4_X1 _24128_ (.A1(_14424_),
    .A2(_14425_),
    .A3(_14426_),
    .A4(_14427_),
    .ZN(_14428_));
 OAI21_X1 _24129_ (.A(_14270_),
    .B1(_14423_),
    .B2(_14079_),
    .ZN(_14429_));
 NAND2_X1 _24130_ (.A1(_14270_),
    .A2(_13981_),
    .ZN(_14430_));
 NAND4_X1 _24131_ (.A1(_14429_),
    .A2(_14272_),
    .A3(_14334_),
    .A4(_14430_),
    .ZN(_14431_));
 INV_X1 _24132_ (.A(_14423_),
    .ZN(_14432_));
 AND2_X1 _24133_ (.A1(_13961_),
    .A2(_14146_),
    .ZN(_14433_));
 INV_X1 _24134_ (.A(_14433_),
    .ZN(_14434_));
 AOI21_X1 _24135_ (.A(_14127_),
    .B1(_14432_),
    .B2(_14434_),
    .ZN(_14435_));
 AND4_X1 _24136_ (.A1(_13997_),
    .A2(_14133_),
    .A3(_14061_),
    .A4(_14278_),
    .ZN(_14436_));
 NOR4_X1 _24137_ (.A1(_14431_),
    .A2(_14435_),
    .A3(_14436_),
    .A4(_14125_),
    .ZN(_14437_));
 NAND4_X1 _24138_ (.A1(_14410_),
    .A2(_14422_),
    .A3(_14428_),
    .A4(_14437_),
    .ZN(_14438_));
 NOR2_X1 _24139_ (.A1(_14402_),
    .A2(_14438_),
    .ZN(_14439_));
 INV_X1 _24140_ (.A(_00992_),
    .ZN(_14440_));
 XNOR2_X1 _24141_ (.A(_14439_),
    .B(_14440_),
    .ZN(_14441_));
 MUX2_X1 _24142_ (.A(_01328_),
    .B(_14441_),
    .S(_14285_),
    .Z(_01083_));
 INV_X1 _24143_ (.A(_14342_),
    .ZN(_14442_));
 AND2_X1 _24144_ (.A1(_14025_),
    .A2(_14041_),
    .ZN(_14443_));
 NOR4_X1 _24145_ (.A1(_14442_),
    .A2(_14443_),
    .A3(_14228_),
    .A4(_14340_),
    .ZN(_14444_));
 AND2_X1 _24146_ (.A1(_14054_),
    .A2(_14055_),
    .ZN(_14445_));
 AOI21_X1 _24147_ (.A(_14065_),
    .B1(_14416_),
    .B2(_14418_),
    .ZN(_14446_));
 AOI211_X1 _24148_ (.A(_14445_),
    .B(_14446_),
    .C1(_14225_),
    .C2(_14141_),
    .ZN(_14447_));
 OAI21_X1 _24149_ (.A(_14067_),
    .B1(_14332_),
    .B2(_14267_),
    .ZN(_14448_));
 AND3_X1 _24150_ (.A1(_14448_),
    .A2(_14071_),
    .A3(_14243_),
    .ZN(_14449_));
 AND2_X1 _24151_ (.A1(_14027_),
    .A2(_14078_),
    .ZN(_14450_));
 AOI211_X1 _24152_ (.A(_14450_),
    .B(_14247_),
    .C1(_14252_),
    .C2(_14141_),
    .ZN(_14451_));
 AND4_X1 _24153_ (.A1(_14444_),
    .A2(_14447_),
    .A3(_14449_),
    .A4(_14451_),
    .ZN(_14452_));
 AOI21_X1 _24154_ (.A(_14116_),
    .B1(_14273_),
    .B2(_14104_),
    .ZN(_14453_));
 OAI21_X1 _24155_ (.A(_14258_),
    .B1(_14177_),
    .B2(_14043_),
    .ZN(_14454_));
 OAI21_X1 _24156_ (.A(_14108_),
    .B1(_13959_),
    .B2(_14236_),
    .ZN(_14455_));
 OAI211_X1 _24157_ (.A(_14454_),
    .B(_14455_),
    .C1(_14119_),
    .C2(_14109_),
    .ZN(_14456_));
 AOI211_X1 _24158_ (.A(_14453_),
    .B(_14456_),
    .C1(_13962_),
    .C2(_14263_),
    .ZN(_14457_));
 OAI211_X1 _24159_ (.A(_14270_),
    .B(_14267_),
    .C1(_14146_),
    .C2(_14100_),
    .ZN(_14458_));
 OAI21_X1 _24160_ (.A(_14270_),
    .B1(_14129_),
    .B2(_14056_),
    .ZN(_14459_));
 AND4_X1 _24161_ (.A1(_14096_),
    .A2(_14458_),
    .A3(_14430_),
    .A4(_14459_),
    .ZN(_14460_));
 AND2_X1 _24162_ (.A1(_14189_),
    .A2(_14087_),
    .ZN(_14461_));
 AND2_X1 _24163_ (.A1(_14215_),
    .A2(_14087_),
    .ZN(_14462_));
 NOR2_X1 _24164_ (.A1(_14461_),
    .A2(_14462_),
    .ZN(_14463_));
 NAND2_X1 _24165_ (.A1(_14133_),
    .A2(_14267_),
    .ZN(_14464_));
 OAI211_X1 _24166_ (.A(_13949_),
    .B(_14086_),
    .C1(_14129_),
    .C2(_14278_),
    .ZN(_14465_));
 AND3_X1 _24167_ (.A1(_14463_),
    .A2(_14464_),
    .A3(_14465_),
    .ZN(_14466_));
 AND4_X1 _24168_ (.A1(_14452_),
    .A2(_14457_),
    .A3(_14460_),
    .A4(_14466_),
    .ZN(_14467_));
 INV_X1 _24169_ (.A(_14182_),
    .ZN(_14468_));
 OAI21_X1 _24170_ (.A(_14143_),
    .B1(_14083_),
    .B2(_14237_),
    .ZN(_14469_));
 OAI21_X1 _24171_ (.A(_14137_),
    .B1(_14095_),
    .B2(_14056_),
    .ZN(_14470_));
 OAI21_X1 _24172_ (.A(_14137_),
    .B1(_14319_),
    .B2(_14237_),
    .ZN(_14471_));
 AND4_X1 _24173_ (.A1(_14468_),
    .A2(_14469_),
    .A3(_14470_),
    .A4(_14471_),
    .ZN(_14472_));
 AOI211_X1 _24174_ (.A(_14294_),
    .B(_14296_),
    .C1(_14237_),
    .C2(_13994_),
    .ZN(_14473_));
 OAI21_X1 _24175_ (.A(_14199_),
    .B1(_14226_),
    .B2(_14118_),
    .ZN(_14474_));
 AND2_X1 _24176_ (.A1(_13967_),
    .A2(_13978_),
    .ZN(_14475_));
 AND2_X1 _24177_ (.A1(_13967_),
    .A2(_14095_),
    .ZN(_14476_));
 AND2_X1 _24178_ (.A1(_13967_),
    .A2(_14118_),
    .ZN(_14477_));
 NOR3_X1 _24179_ (.A1(_14475_),
    .A2(_14476_),
    .A3(_14477_),
    .ZN(_14478_));
 AND4_X1 _24180_ (.A1(_14293_),
    .A2(_14473_),
    .A3(_14474_),
    .A4(_14478_),
    .ZN(_14479_));
 NAND2_X1 _24181_ (.A1(_14171_),
    .A2(_14423_),
    .ZN(_14480_));
 OAI21_X1 _24182_ (.A(_14171_),
    .B1(_14177_),
    .B2(_13978_),
    .ZN(_14481_));
 OAI211_X1 _24183_ (.A(_14480_),
    .B(_14481_),
    .C1(_14185_),
    .C2(_14324_),
    .ZN(_14482_));
 AND4_X1 _24184_ (.A1(_13971_),
    .A2(_14022_),
    .A3(_14004_),
    .A4(_14136_),
    .ZN(_14483_));
 OR2_X1 _24185_ (.A1(_14176_),
    .A2(_14483_),
    .ZN(_14484_));
 NOR4_X1 _24186_ (.A1(_14482_),
    .A2(_14484_),
    .A3(_14152_),
    .A4(_14375_),
    .ZN(_14485_));
 NAND2_X1 _24187_ (.A1(_14246_),
    .A2(_13952_),
    .ZN(_14486_));
 OAI221_X1 _24188_ (.A(_14486_),
    .B1(_14312_),
    .B2(_14191_),
    .C1(_14220_),
    .C2(_11040_),
    .ZN(_14487_));
 AOI21_X1 _24189_ (.A(_14010_),
    .B1(_14420_),
    .B2(_14034_),
    .ZN(_14488_));
 NOR4_X1 _24190_ (.A1(_14487_),
    .A2(_14488_),
    .A3(_14016_),
    .A4(_14217_),
    .ZN(_14489_));
 AND4_X1 _24191_ (.A1(_14472_),
    .A2(_14479_),
    .A3(_14485_),
    .A4(_14489_),
    .ZN(_14490_));
 AND3_X1 _24192_ (.A1(_14467_),
    .A2(_00993_),
    .A3(_14490_),
    .ZN(_14491_));
 AOI21_X1 _24193_ (.A(_00993_),
    .B1(_14467_),
    .B2(_14490_),
    .ZN(_14492_));
 NOR2_X1 _24194_ (.A1(_14491_),
    .A2(_14492_),
    .ZN(_14493_));
 MUX2_X1 _24195_ (.A(_01203_),
    .B(_14493_),
    .S(_14285_),
    .Z(_01084_));
 AOI21_X1 _24196_ (.A(_14130_),
    .B1(_14187_),
    .B2(_14179_),
    .ZN(_14494_));
 AOI21_X1 _24197_ (.A(_14494_),
    .B1(_14252_),
    .B2(_13978_),
    .ZN(_14495_));
 AOI22_X1 _24198_ (.A1(_14301_),
    .A2(_14146_),
    .B1(_13953_),
    .B2(_14215_),
    .ZN(_14496_));
 NAND4_X1 _24199_ (.A1(_14495_),
    .A2(_14496_),
    .A3(_14090_),
    .A4(_14342_),
    .ZN(_14497_));
 INV_X1 _24200_ (.A(_14168_),
    .ZN(_14498_));
 NAND3_X1 _24201_ (.A1(_14236_),
    .A2(_13949_),
    .A3(_14145_),
    .ZN(_14499_));
 AND2_X1 _24202_ (.A1(_14498_),
    .A2(_14499_),
    .ZN(_14500_));
 OAI21_X1 _24203_ (.A(_14263_),
    .B1(_13978_),
    .B2(_14132_),
    .ZN(_14501_));
 NOR2_X1 _24204_ (.A1(_14318_),
    .A2(_13973_),
    .ZN(_14502_));
 OAI21_X1 _24205_ (.A(_14143_),
    .B1(_14502_),
    .B2(_14246_),
    .ZN(_14503_));
 OAI21_X1 _24206_ (.A(_14250_),
    .B1(_14417_),
    .B2(_13962_),
    .ZN(_14504_));
 NAND4_X1 _24207_ (.A1(_14500_),
    .A2(_14501_),
    .A3(_14503_),
    .A4(_14504_),
    .ZN(_14505_));
 OAI211_X1 _24208_ (.A(_14272_),
    .B(_14241_),
    .C1(_14356_),
    .C2(_14113_),
    .ZN(_14506_));
 AND2_X1 _24209_ (.A1(_14092_),
    .A2(_13952_),
    .ZN(_14507_));
 OR2_X1 _24210_ (.A1(_14507_),
    .A2(_14404_),
    .ZN(_14508_));
 NOR4_X1 _24211_ (.A1(_14497_),
    .A2(_14505_),
    .A3(_14506_),
    .A4(_14508_),
    .ZN(_14509_));
 OAI21_X1 _24212_ (.A(_14199_),
    .B1(_13978_),
    .B2(_14056_),
    .ZN(_14510_));
 NAND4_X1 _24213_ (.A1(_14199_),
    .A2(_13997_),
    .A3(_14061_),
    .A4(_14278_),
    .ZN(_14511_));
 OAI211_X1 _24214_ (.A(_14510_),
    .B(_14511_),
    .C1(_13990_),
    .C2(_14119_),
    .ZN(_14512_));
 AOI21_X1 _24215_ (.A(_13990_),
    .B1(_14432_),
    .B2(_14434_),
    .ZN(_14513_));
 NOR3_X1 _24216_ (.A1(_14512_),
    .A2(_14123_),
    .A3(_14513_),
    .ZN(_14514_));
 NAND2_X1 _24217_ (.A1(_14252_),
    .A2(_14079_),
    .ZN(_14515_));
 OAI221_X1 _24218_ (.A(_14515_),
    .B1(_14112_),
    .B2(_14127_),
    .C1(_14119_),
    .C2(_13968_),
    .ZN(_14516_));
 AND2_X1 _24219_ (.A1(_14141_),
    .A2(_14054_),
    .ZN(_14517_));
 AND2_X1 _24220_ (.A1(_14517_),
    .A2(_14007_),
    .ZN(_14518_));
 AND3_X1 _24221_ (.A1(_14083_),
    .A2(_14225_),
    .A3(_14061_),
    .ZN(_14519_));
 NOR4_X1 _24222_ (.A1(_14516_),
    .A2(_14484_),
    .A3(_14518_),
    .A4(_14519_),
    .ZN(_14520_));
 AND2_X1 _24223_ (.A1(_14054_),
    .A2(_14236_),
    .ZN(_14521_));
 INV_X1 _24224_ (.A(_14521_),
    .ZN(_14522_));
 NAND3_X1 _24225_ (.A1(_14077_),
    .A2(_14026_),
    .A3(_13983_),
    .ZN(_14523_));
 AND3_X1 _24226_ (.A1(_14522_),
    .A2(_14220_),
    .A3(_14523_),
    .ZN(_14524_));
 NAND2_X1 _24227_ (.A1(_14171_),
    .A2(_14092_),
    .ZN(_14525_));
 NAND2_X1 _24228_ (.A1(_14525_),
    .A2(_14126_),
    .ZN(_14526_));
 AND2_X1 _24229_ (.A1(_14054_),
    .A2(_14025_),
    .ZN(_14527_));
 NOR4_X1 _24230_ (.A1(_14156_),
    .A2(_14526_),
    .A3(_14389_),
    .A4(_14527_),
    .ZN(_14528_));
 AOI22_X1 _24231_ (.A1(_13994_),
    .A2(_14189_),
    .B1(_13988_),
    .B2(_14252_),
    .ZN(_14529_));
 AOI22_X1 _24232_ (.A1(_14013_),
    .A2(_14137_),
    .B1(_14189_),
    .B2(_14133_),
    .ZN(_14530_));
 AND4_X1 _24233_ (.A1(_14524_),
    .A2(_14528_),
    .A3(_14529_),
    .A4(_14530_),
    .ZN(_14531_));
 NAND4_X1 _24234_ (.A1(_14509_),
    .A2(_14514_),
    .A3(_14520_),
    .A4(_14531_),
    .ZN(_14532_));
 AOI211_X1 _24235_ (.A(_14003_),
    .B(_14179_),
    .C1(_14140_),
    .C2(_13995_),
    .ZN(_14533_));
 AOI211_X1 _24236_ (.A(_14021_),
    .B(_14533_),
    .C1(_14018_),
    .C2(_14317_),
    .ZN(_14534_));
 OAI21_X1 _24237_ (.A(_14096_),
    .B1(_14065_),
    .B2(_14104_),
    .ZN(_14535_));
 NOR2_X1 _24238_ (.A1(_14535_),
    .A2(_14443_),
    .ZN(_14536_));
 AOI22_X1 _24239_ (.A1(_14025_),
    .A2(_14171_),
    .B1(_14143_),
    .B2(_14056_),
    .ZN(_14537_));
 OAI21_X1 _24240_ (.A(_14059_),
    .B1(_14160_),
    .B2(_14252_),
    .ZN(_14538_));
 NAND4_X1 _24241_ (.A1(_14534_),
    .A2(_14536_),
    .A3(_14537_),
    .A4(_14538_),
    .ZN(_14539_));
 AOI22_X1 _24242_ (.A1(_14022_),
    .A2(_13994_),
    .B1(_14143_),
    .B2(_14236_),
    .ZN(_14540_));
 OAI211_X1 _24243_ (.A(_14430_),
    .B(_14540_),
    .C1(_14185_),
    .C2(_14187_),
    .ZN(_14541_));
 AND2_X1 _24244_ (.A1(_14006_),
    .A2(_14118_),
    .ZN(_14542_));
 NOR2_X1 _24245_ (.A1(_14169_),
    .A2(_14542_),
    .ZN(_14543_));
 NAND2_X1 _24246_ (.A1(_13953_),
    .A2(_14417_),
    .ZN(_14544_));
 OAI21_X1 _24247_ (.A(_14317_),
    .B1(_13959_),
    .B2(_14059_),
    .ZN(_14545_));
 AOI22_X1 _24248_ (.A1(_14160_),
    .A2(_14079_),
    .B1(_14091_),
    .B2(_14015_),
    .ZN(_14546_));
 NAND4_X1 _24249_ (.A1(_14543_),
    .A2(_14544_),
    .A3(_14545_),
    .A4(_14546_),
    .ZN(_14547_));
 AND3_X1 _24250_ (.A1(_14095_),
    .A2(_13965_),
    .A3(_14086_),
    .ZN(_14548_));
 AND2_X1 _24251_ (.A1(_14108_),
    .A2(_14055_),
    .ZN(_14549_));
 AOI211_X1 _24252_ (.A(_14548_),
    .B(_14549_),
    .C1(_14013_),
    .C2(_14258_),
    .ZN(_14550_));
 OAI21_X1 _24253_ (.A(_14258_),
    .B1(_14025_),
    .B2(_14237_),
    .ZN(_14551_));
 OAI211_X1 _24254_ (.A(_14550_),
    .B(_14551_),
    .C1(_14049_),
    .C2(_14130_),
    .ZN(_14552_));
 OR4_X1 _24255_ (.A1(_14539_),
    .A2(_14541_),
    .A3(_14547_),
    .A4(_14552_),
    .ZN(_14553_));
 NOR2_X1 _24256_ (.A1(_14532_),
    .A2(_14553_),
    .ZN(_14554_));
 XOR2_X1 _24257_ (.A(_14554_),
    .B(_00994_),
    .Z(_14555_));
 MUX2_X1 _24258_ (.A(_01204_),
    .B(_14555_),
    .S(_14285_),
    .Z(_01085_));
 AOI211_X1 _24259_ (.A(_14161_),
    .B(_14375_),
    .C1(_14160_),
    .C2(_14129_),
    .ZN(_14556_));
 NAND2_X1 _24260_ (.A1(_14160_),
    .A2(_14079_),
    .ZN(_14557_));
 OAI211_X1 _24261_ (.A(_14556_),
    .B(_14557_),
    .C1(_14179_),
    .C2(_14101_),
    .ZN(_14558_));
 OAI21_X1 _24262_ (.A(_14143_),
    .B1(_14200_),
    .B2(_14226_),
    .ZN(_14559_));
 OAI211_X1 _24263_ (.A(_13983_),
    .B(_14145_),
    .C1(_14031_),
    .C2(_13988_),
    .ZN(_14560_));
 OAI211_X1 _24264_ (.A(_14559_),
    .B(_14560_),
    .C1(_14434_),
    .C2(_14183_),
    .ZN(_14561_));
 OAI211_X1 _24265_ (.A(_14194_),
    .B(_14145_),
    .C1(_14129_),
    .C2(_14022_),
    .ZN(_14562_));
 OAI211_X1 _24266_ (.A(_14562_),
    .B(_14190_),
    .C1(_14187_),
    .C2(_14318_),
    .ZN(_14563_));
 OAI211_X1 _24267_ (.A(_14171_),
    .B(_17086_),
    .C1(_14100_),
    .C2(_13969_),
    .ZN(_14564_));
 OAI211_X1 _24268_ (.A(_13949_),
    .B(_14145_),
    .C1(_14056_),
    .C2(_14118_),
    .ZN(_14565_));
 OAI211_X1 _24269_ (.A(_14564_),
    .B(_14565_),
    .C1(_14064_),
    .C2(_14324_),
    .ZN(_14566_));
 NOR4_X1 _24270_ (.A1(_14558_),
    .A2(_14561_),
    .A3(_14563_),
    .A4(_14566_),
    .ZN(_14567_));
 OR3_X1 _24271_ (.A1(_14042_),
    .A2(_14044_),
    .A3(_14228_),
    .ZN(_14568_));
 NOR3_X1 _24272_ (.A1(_14568_),
    .A2(_14442_),
    .A3(_14341_),
    .ZN(_14569_));
 NAND3_X1 _24273_ (.A1(_14092_),
    .A2(_14026_),
    .A3(_14194_),
    .ZN(_14570_));
 OAI211_X1 _24274_ (.A(_14348_),
    .B(_14570_),
    .C1(_14065_),
    .C2(_14097_),
    .ZN(_14571_));
 NAND2_X1 _24275_ (.A1(_14054_),
    .A2(_14246_),
    .ZN(_14572_));
 NAND2_X1 _24276_ (.A1(_14054_),
    .A2(_14031_),
    .ZN(_14573_));
 OAI211_X1 _24277_ (.A(_14572_),
    .B(_14573_),
    .C1(_14065_),
    .C2(_14244_),
    .ZN(_14574_));
 AOI211_X1 _24278_ (.A(_14571_),
    .B(_14574_),
    .C1(_14225_),
    .C2(_14155_),
    .ZN(_14575_));
 NAND2_X1 _24279_ (.A1(_14020_),
    .A2(_14250_),
    .ZN(_14576_));
 OAI21_X1 _24280_ (.A(_14250_),
    .B1(_14423_),
    .B2(_14076_),
    .ZN(_14577_));
 NAND2_X1 _24281_ (.A1(_14250_),
    .A2(_14237_),
    .ZN(_14578_));
 AND4_X1 _24282_ (.A1(_14576_),
    .A2(_14577_),
    .A3(_14578_),
    .A4(_14355_),
    .ZN(_14579_));
 OAI21_X1 _24283_ (.A(_14427_),
    .B1(_14032_),
    .B2(_14029_),
    .ZN(_14580_));
 AND2_X1 _24284_ (.A1(_14252_),
    .A2(_14265_),
    .ZN(_14581_));
 NOR3_X1 _24285_ (.A1(_14580_),
    .A2(_14248_),
    .A3(_14581_),
    .ZN(_14582_));
 AND4_X1 _24286_ (.A1(_14569_),
    .A2(_14575_),
    .A3(_14579_),
    .A4(_14582_),
    .ZN(_14583_));
 AOI21_X1 _24287_ (.A(_14116_),
    .B1(_14432_),
    .B2(_14434_),
    .ZN(_14584_));
 AOI21_X1 _24288_ (.A(_14584_),
    .B1(_14063_),
    .B2(_14263_),
    .ZN(_14585_));
 OR2_X1 _24289_ (.A1(_14109_),
    .A2(_14113_),
    .ZN(_14586_));
 NAND2_X1 _24290_ (.A1(_14258_),
    .A2(_14132_),
    .ZN(_14587_));
 AND4_X1 _24291_ (.A1(_14586_),
    .A2(_14257_),
    .A3(_14587_),
    .A4(_14411_),
    .ZN(_14588_));
 AOI21_X1 _24292_ (.A(_14098_),
    .B1(_14119_),
    .B2(_14104_),
    .ZN(_14589_));
 AND2_X1 _24293_ (.A1(_14270_),
    .A2(_14013_),
    .ZN(_14590_));
 AND2_X1 _24294_ (.A1(_14091_),
    .A2(_14076_),
    .ZN(_14591_));
 NOR4_X1 _24295_ (.A1(_14589_),
    .A2(_14102_),
    .A3(_14590_),
    .A4(_14591_),
    .ZN(_14592_));
 OAI21_X1 _24296_ (.A(_14133_),
    .B1(_14092_),
    .B2(_14172_),
    .ZN(_14593_));
 INV_X1 _24297_ (.A(_14462_),
    .ZN(_14594_));
 AND3_X1 _24298_ (.A1(_14593_),
    .A2(_14277_),
    .A3(_14594_),
    .ZN(_14595_));
 AND4_X1 _24299_ (.A1(_14585_),
    .A2(_14588_),
    .A3(_14592_),
    .A4(_14595_),
    .ZN(_14596_));
 OAI21_X1 _24300_ (.A(_13994_),
    .B1(_14200_),
    .B2(_14226_),
    .ZN(_14597_));
 AND2_X1 _24301_ (.A1(_14189_),
    .A2(_14198_),
    .ZN(_14598_));
 AOI211_X1 _24302_ (.A(_14204_),
    .B(_14598_),
    .C1(_14199_),
    .C2(_14215_),
    .ZN(_14599_));
 OAI21_X1 _24303_ (.A(_14199_),
    .B1(_14092_),
    .B2(_14020_),
    .ZN(_14600_));
 AND2_X1 _24304_ (.A1(_14599_),
    .A2(_14600_),
    .ZN(_14601_));
 OAI21_X1 _24305_ (.A(_13994_),
    .B1(_14423_),
    .B2(_14433_),
    .ZN(_14602_));
 OAI21_X1 _24306_ (.A(_13953_),
    .B1(_14423_),
    .B2(_14025_),
    .ZN(_14603_));
 OAI21_X1 _24307_ (.A(_14317_),
    .B1(_14319_),
    .B2(_14059_),
    .ZN(_14604_));
 OAI21_X1 _24308_ (.A(_14317_),
    .B1(_14013_),
    .B2(_14118_),
    .ZN(_14605_));
 OAI211_X1 _24309_ (.A(_13952_),
    .B(_14278_),
    .C1(_11040_),
    .C2(_11046_),
    .ZN(_14606_));
 AND4_X1 _24310_ (.A1(_14603_),
    .A2(_14604_),
    .A3(_14605_),
    .A4(_14606_),
    .ZN(_14607_));
 AND4_X1 _24311_ (.A1(_14597_),
    .A2(_14601_),
    .A3(_14602_),
    .A4(_14607_),
    .ZN(_14608_));
 NAND4_X1 _24312_ (.A1(_14567_),
    .A2(_14583_),
    .A3(_14596_),
    .A4(_14608_),
    .ZN(_14609_));
 NOR2_X1 _24313_ (.A1(_14609_),
    .A2(_14164_),
    .ZN(_14610_));
 XOR2_X1 _24314_ (.A(_14610_),
    .B(_00995_),
    .Z(_14611_));
 MUX2_X1 _24315_ (.A(_01205_),
    .B(_14611_),
    .S(_14285_),
    .Z(_01086_));
 AND2_X1 _24316_ (.A1(_14091_),
    .A2(_14246_),
    .ZN(_14612_));
 NAND2_X1 _24317_ (.A1(_14091_),
    .A2(_14022_),
    .ZN(_14613_));
 OAI211_X1 _24318_ (.A(_14094_),
    .B(_14613_),
    .C1(_14098_),
    .C2(_14119_),
    .ZN(_14614_));
 AOI211_X1 _24319_ (.A(_14612_),
    .B(_14614_),
    .C1(_14079_),
    .C2(_14270_),
    .ZN(_14615_));
 OAI211_X1 _24320_ (.A(_14133_),
    .B(_14278_),
    .C1(_11040_),
    .C2(_14100_),
    .ZN(_14616_));
 AND2_X1 _24321_ (.A1(_14616_),
    .A2(_14275_),
    .ZN(_14617_));
 AND4_X1 _24322_ (.A1(_14277_),
    .A2(_14615_),
    .A3(_14463_),
    .A4(_14617_),
    .ZN(_14618_));
 NAND4_X1 _24323_ (.A1(_14522_),
    .A2(_14345_),
    .A3(_14346_),
    .A4(_14573_),
    .ZN(_14619_));
 NAND3_X1 _24324_ (.A1(_14141_),
    .A2(_14047_),
    .A3(_14007_),
    .ZN(_14620_));
 OAI211_X1 _24325_ (.A(_14620_),
    .B(_14234_),
    .C1(_14049_),
    .C2(_14244_),
    .ZN(_14621_));
 AOI21_X1 _24326_ (.A(_14065_),
    .B1(_14119_),
    .B2(_13979_),
    .ZN(_14622_));
 NOR4_X1 _24327_ (.A1(_14619_),
    .A2(_14518_),
    .A3(_14621_),
    .A4(_14622_),
    .ZN(_14623_));
 NAND4_X1 _24328_ (.A1(_14071_),
    .A2(_14074_),
    .A3(_14355_),
    .A4(_14424_),
    .ZN(_14624_));
 AND3_X1 _24329_ (.A1(_14252_),
    .A2(_11040_),
    .A3(_14278_),
    .ZN(_14625_));
 AOI21_X1 _24330_ (.A(_14029_),
    .B1(_14418_),
    .B2(_14412_),
    .ZN(_14626_));
 NOR4_X1 _24331_ (.A1(_14624_),
    .A2(_14625_),
    .A3(_14581_),
    .A4(_14626_),
    .ZN(_14627_));
 AND4_X1 _24332_ (.A1(_11039_),
    .A2(_14194_),
    .A3(_14086_),
    .A4(_14008_),
    .ZN(_14628_));
 AOI211_X1 _24333_ (.A(_14628_),
    .B(_14548_),
    .C1(_14177_),
    .C2(_14258_),
    .ZN(_14629_));
 OAI21_X1 _24334_ (.A(_14258_),
    .B1(_14184_),
    .B2(_14031_),
    .ZN(_14630_));
 OAI21_X1 _24335_ (.A(_14263_),
    .B1(_14092_),
    .B2(_14020_),
    .ZN(_14631_));
 OAI21_X1 _24336_ (.A(_14263_),
    .B1(_14015_),
    .B2(_14237_),
    .ZN(_14632_));
 AND4_X1 _24337_ (.A1(_14629_),
    .A2(_14630_),
    .A3(_14631_),
    .A4(_14632_),
    .ZN(_14633_));
 NAND4_X1 _24338_ (.A1(_14618_),
    .A2(_14623_),
    .A3(_14627_),
    .A4(_14633_),
    .ZN(_14634_));
 AND2_X1 _24339_ (.A1(_14177_),
    .A2(_14317_),
    .ZN(_14635_));
 AND2_X1 _24340_ (.A1(_13978_),
    .A2(_14006_),
    .ZN(_14636_));
 OR4_X1 _24341_ (.A1(_14635_),
    .A2(_14310_),
    .A3(_14636_),
    .A4(_14542_),
    .ZN(_14637_));
 NAND2_X1 _24342_ (.A1(_14069_),
    .A2(_13953_),
    .ZN(_14638_));
 NAND4_X1 _24343_ (.A1(_14486_),
    .A2(_14220_),
    .A3(_14638_),
    .A4(_14544_),
    .ZN(_14639_));
 NOR4_X1 _24344_ (.A1(_14637_),
    .A2(_14639_),
    .A3(_14214_),
    .A4(_14012_),
    .ZN(_14640_));
 NOR2_X1 _24345_ (.A1(_14475_),
    .A2(_14476_),
    .ZN(_14641_));
 OAI211_X1 _24346_ (.A(_14194_),
    .B(_13950_),
    .C1(_14031_),
    .C2(_13988_),
    .ZN(_14642_));
 OAI211_X1 _24347_ (.A(_14641_),
    .B(_14642_),
    .C1(_14314_),
    .C2(_13968_),
    .ZN(_14643_));
 NAND3_X1 _24348_ (.A1(_14199_),
    .A2(_14278_),
    .A3(_13973_),
    .ZN(_14644_));
 NAND2_X1 _24349_ (.A1(_14199_),
    .A2(_14129_),
    .ZN(_14645_));
 OAI211_X1 _24350_ (.A(_14644_),
    .B(_14645_),
    .C1(_14112_),
    .C2(_13990_),
    .ZN(_14646_));
 AOI211_X1 _24351_ (.A(_14191_),
    .B(_13990_),
    .C1(_14146_),
    .C2(_14100_),
    .ZN(_14647_));
 NOR4_X1 _24352_ (.A1(_14643_),
    .A2(_14598_),
    .A3(_14646_),
    .A4(_14647_),
    .ZN(_14648_));
 NAND3_X1 _24353_ (.A1(_14189_),
    .A2(_13983_),
    .A3(_14145_),
    .ZN(_14649_));
 OAI21_X1 _24354_ (.A(_14137_),
    .B1(_14184_),
    .B2(_14502_),
    .ZN(_14650_));
 OAI211_X1 _24355_ (.A(_14194_),
    .B(_14145_),
    .C1(_14043_),
    .C2(_14265_),
    .ZN(_14651_));
 OAI21_X1 _24356_ (.A(_14143_),
    .B1(_14200_),
    .B2(_14177_),
    .ZN(_14652_));
 AND4_X1 _24357_ (.A1(_14649_),
    .A2(_14650_),
    .A3(_14651_),
    .A4(_14652_),
    .ZN(_14653_));
 NAND2_X1 _24358_ (.A1(_14160_),
    .A2(_14129_),
    .ZN(_14654_));
 OAI221_X1 _24359_ (.A(_14160_),
    .B1(_14146_),
    .B2(_14100_),
    .C1(_14267_),
    .C2(_13962_),
    .ZN(_14655_));
 OAI21_X1 _24360_ (.A(_14171_),
    .B1(_14141_),
    .B2(_14118_),
    .ZN(_14656_));
 AND4_X1 _24361_ (.A1(_14500_),
    .A2(_14654_),
    .A3(_14655_),
    .A4(_14656_),
    .ZN(_14657_));
 NAND4_X1 _24362_ (.A1(_14640_),
    .A2(_14648_),
    .A3(_14653_),
    .A4(_14657_),
    .ZN(_14658_));
 NOR2_X1 _24363_ (.A1(_14634_),
    .A2(_14658_),
    .ZN(_14659_));
 XOR2_X1 _24364_ (.A(_14659_),
    .B(_00996_),
    .Z(_14660_));
 MUX2_X1 _24365_ (.A(_01206_),
    .B(_14660_),
    .S(_14285_),
    .Z(_01087_));
 INV_X1 _24366_ (.A(_17096_),
    .ZN(_14661_));
 AND2_X1 _24367_ (.A1(_14661_),
    .A2(_17095_),
    .ZN(_14662_));
 INV_X1 _24368_ (.A(_17094_),
    .ZN(_14663_));
 AND2_X1 _24369_ (.A1(_14663_),
    .A2(_17093_),
    .ZN(_14664_));
 CLKBUF_X2 _24370_ (.A(_14664_),
    .Z(_14665_));
 AND2_X1 _24371_ (.A1(_14662_),
    .A2(_14665_),
    .ZN(_14666_));
 INV_X2 _24372_ (.A(_14666_),
    .ZN(_14667_));
 INV_X1 _24373_ (.A(_17089_),
    .ZN(_14668_));
 NOR2_X1 _24374_ (.A1(_14668_),
    .A2(_17092_),
    .ZN(_14669_));
 AND2_X1 _24375_ (.A1(_14669_),
    .A2(_17078_),
    .ZN(_14670_));
 BUF_X2 _24376_ (.A(_14670_),
    .Z(_14671_));
 INV_X1 _24377_ (.A(_14671_),
    .ZN(_14672_));
 NOR2_X2 _24378_ (.A1(_17093_),
    .A2(_17094_),
    .ZN(_14673_));
 AND2_X1 _24379_ (.A1(_14662_),
    .A2(_14673_),
    .ZN(_14674_));
 BUF_X2 _24380_ (.A(_14674_),
    .Z(_14675_));
 INV_X2 _24381_ (.A(_14675_),
    .ZN(_14676_));
 NOR2_X2 _24382_ (.A1(_17089_),
    .A2(_17092_),
    .ZN(_14677_));
 AND2_X2 _24383_ (.A1(_14677_),
    .A2(_09451_),
    .ZN(_14678_));
 INV_X1 _24384_ (.A(_14678_),
    .ZN(_14679_));
 OAI22_X1 _24385_ (.A1(_14667_),
    .A2(_14672_),
    .B1(_14676_),
    .B2(_14679_),
    .ZN(_14680_));
 AND2_X2 _24386_ (.A1(_14669_),
    .A2(_09451_),
    .ZN(_14681_));
 NOR2_X1 _24387_ (.A1(_14663_),
    .A2(_17093_),
    .ZN(_14682_));
 AND2_X1 _24388_ (.A1(_14662_),
    .A2(_14682_),
    .ZN(_14683_));
 CLKBUF_X2 _24389_ (.A(_14683_),
    .Z(_14684_));
 AND2_X1 _24390_ (.A1(_17089_),
    .A2(_17092_),
    .ZN(_14685_));
 AND2_X1 _24391_ (.A1(_14685_),
    .A2(_09451_),
    .ZN(_14686_));
 BUF_X2 _24392_ (.A(_14686_),
    .Z(_14687_));
 AND2_X1 _24393_ (.A1(_17093_),
    .A2(_17094_),
    .ZN(_14688_));
 NOR2_X1 _24394_ (.A1(_17095_),
    .A2(_17096_),
    .ZN(_14689_));
 AND2_X2 _24395_ (.A1(_14688_),
    .A2(_14689_),
    .ZN(_14690_));
 BUF_X2 _24396_ (.A(_14690_),
    .Z(_14691_));
 AOI221_X4 _24397_ (.A(_14680_),
    .B1(_14681_),
    .B2(_14684_),
    .C1(_14687_),
    .C2(_14691_),
    .ZN(_14692_));
 AND2_X1 _24398_ (.A1(_17095_),
    .A2(_17096_),
    .ZN(_14693_));
 CLKBUF_X2 _24399_ (.A(_14693_),
    .Z(_14694_));
 AND2_X1 _24400_ (.A1(_14694_),
    .A2(_14673_),
    .ZN(_14695_));
 AND2_X1 _24401_ (.A1(_14686_),
    .A2(_14695_),
    .ZN(_14696_));
 AND2_X1 _24402_ (.A1(_14664_),
    .A2(_14693_),
    .ZN(_14697_));
 CLKBUF_X2 _24403_ (.A(_14697_),
    .Z(_14698_));
 INV_X1 _24404_ (.A(_17092_),
    .ZN(_14699_));
 NOR2_X2 _24405_ (.A1(_14699_),
    .A2(_17089_),
    .ZN(_14700_));
 CLKBUF_X2 _24406_ (.A(_14700_),
    .Z(_14701_));
 AND2_X1 _24407_ (.A1(_14700_),
    .A2(_17067_),
    .ZN(_14702_));
 CLKBUF_X2 _24408_ (.A(_14695_),
    .Z(_14703_));
 AOI221_X4 _24409_ (.A(_14696_),
    .B1(_14698_),
    .B2(_14701_),
    .C1(_14702_),
    .C2(_14703_),
    .ZN(_14704_));
 AND2_X2 _24410_ (.A1(_14689_),
    .A2(_14673_),
    .ZN(_14705_));
 BUF_X2 _24411_ (.A(_14705_),
    .Z(_14706_));
 NOR2_X2 _24412_ (.A1(_17067_),
    .A2(_17078_),
    .ZN(_14707_));
 INV_X1 _24413_ (.A(_14707_),
    .ZN(_14708_));
 CLKBUF_X2 _24414_ (.A(_14685_),
    .Z(_14709_));
 NAND2_X1 _24415_ (.A1(_14708_),
    .A2(_14709_),
    .ZN(_14710_));
 AND2_X1 _24416_ (.A1(_17067_),
    .A2(_17078_),
    .ZN(_14711_));
 BUF_X2 _24417_ (.A(_14711_),
    .Z(_14712_));
 NOR2_X1 _24418_ (.A1(_14710_),
    .A2(_14712_),
    .ZN(_14713_));
 AND2_X1 _24419_ (.A1(_14700_),
    .A2(_17078_),
    .ZN(_14714_));
 OAI21_X1 _24420_ (.A(_14706_),
    .B1(_14713_),
    .B2(_14714_),
    .ZN(_14715_));
 AND2_X2 _24421_ (.A1(_14662_),
    .A2(_14688_),
    .ZN(_14716_));
 BUF_X2 _24422_ (.A(_14716_),
    .Z(_14717_));
 BUF_X2 _24423_ (.A(_14669_),
    .Z(_14718_));
 AND2_X2 _24424_ (.A1(_14718_),
    .A2(_17067_),
    .ZN(_14719_));
 AND2_X1 _24425_ (.A1(_14677_),
    .A2(_17067_),
    .ZN(_14720_));
 OAI21_X1 _24426_ (.A(_14717_),
    .B1(_14719_),
    .B2(_14720_),
    .ZN(_14721_));
 AND4_X1 _24427_ (.A1(_14692_),
    .A2(_14704_),
    .A3(_14715_),
    .A4(_14721_),
    .ZN(_14722_));
 NOR2_X1 _24428_ (.A1(_14661_),
    .A2(_17095_),
    .ZN(_14723_));
 AND2_X1 _24429_ (.A1(_14664_),
    .A2(_14723_),
    .ZN(_14724_));
 CLKBUF_X2 _24430_ (.A(_14724_),
    .Z(_14725_));
 INV_X1 _24431_ (.A(_14677_),
    .ZN(_14726_));
 NOR2_X1 _24432_ (.A1(_14726_),
    .A2(_14712_),
    .ZN(_14727_));
 AND3_X1 _24433_ (.A1(_14725_),
    .A2(_14708_),
    .A3(_14727_),
    .ZN(_14728_));
 AND2_X1 _24434_ (.A1(_14664_),
    .A2(_14689_),
    .ZN(_14729_));
 INV_X2 _24435_ (.A(_14729_),
    .ZN(_14730_));
 NOR2_X1 _24436_ (.A1(_09451_),
    .A2(_17067_),
    .ZN(_14731_));
 CLKBUF_X2 _24437_ (.A(_14731_),
    .Z(_14732_));
 NOR3_X1 _24438_ (.A1(_14732_),
    .A2(_17089_),
    .A3(_14699_),
    .ZN(_14733_));
 INV_X1 _24439_ (.A(_17067_),
    .ZN(_14734_));
 NOR2_X2 _24440_ (.A1(_14734_),
    .A2(_17078_),
    .ZN(_14735_));
 INV_X1 _24441_ (.A(_14735_),
    .ZN(_14736_));
 AND2_X1 _24442_ (.A1(_14733_),
    .A2(_14736_),
    .ZN(_14737_));
 INV_X1 _24443_ (.A(_14737_),
    .ZN(_14738_));
 INV_X2 _24444_ (.A(_14712_),
    .ZN(_14739_));
 NAND2_X2 _24445_ (.A1(_14739_),
    .A2(_14718_),
    .ZN(_14740_));
 NOR2_X1 _24446_ (.A1(_14740_),
    .A2(_14707_),
    .ZN(_14741_));
 INV_X1 _24447_ (.A(_14741_),
    .ZN(_14742_));
 AOI21_X1 _24448_ (.A(_14730_),
    .B1(_14738_),
    .B2(_14742_),
    .ZN(_14743_));
 AND2_X1 _24449_ (.A1(_14685_),
    .A2(_17078_),
    .ZN(_14744_));
 CLKBUF_X2 _24450_ (.A(_14744_),
    .Z(_14745_));
 AOI211_X1 _24451_ (.A(_14728_),
    .B(_14743_),
    .C1(_14745_),
    .C2(_14725_),
    .ZN(_14746_));
 AND2_X1 _24452_ (.A1(_14685_),
    .A2(_14707_),
    .ZN(_14747_));
 BUF_X2 _24453_ (.A(_14747_),
    .Z(_14748_));
 CLKBUF_X2 _24454_ (.A(_14682_),
    .Z(_14749_));
 AND2_X1 _24455_ (.A1(_14749_),
    .A2(_14689_),
    .ZN(_14750_));
 BUF_X2 _24456_ (.A(_14750_),
    .Z(_14751_));
 AND2_X1 _24457_ (.A1(_14709_),
    .A2(_14712_),
    .ZN(_14752_));
 BUF_X2 _24458_ (.A(_14752_),
    .Z(_14753_));
 AOI22_X1 _24459_ (.A1(_14748_),
    .A2(_14751_),
    .B1(_14753_),
    .B2(_14691_),
    .ZN(_14754_));
 AND2_X2 _24460_ (.A1(_14669_),
    .A2(_14707_),
    .ZN(_14755_));
 INV_X1 _24461_ (.A(_14755_),
    .ZN(_14756_));
 INV_X1 _24462_ (.A(_14683_),
    .ZN(_14757_));
 OAI221_X1 _24463_ (.A(_14754_),
    .B1(_14676_),
    .B2(_14756_),
    .C1(_14672_),
    .C2(_14757_),
    .ZN(_14758_));
 AND2_X1 _24464_ (.A1(_14718_),
    .A2(_14735_),
    .ZN(_14759_));
 BUF_X2 _24465_ (.A(_14759_),
    .Z(_14760_));
 AND2_X2 _24466_ (.A1(_14735_),
    .A2(_14700_),
    .ZN(_14761_));
 OAI21_X1 _24467_ (.A(_14706_),
    .B1(_14760_),
    .B2(_14761_),
    .ZN(_14762_));
 AND2_X2 _24468_ (.A1(_14677_),
    .A2(_17078_),
    .ZN(_14763_));
 BUF_X2 _24469_ (.A(_14689_),
    .Z(_14764_));
 NAND3_X1 _24470_ (.A1(_14763_),
    .A2(_14663_),
    .A3(_14764_),
    .ZN(_14765_));
 INV_X1 _24471_ (.A(_14705_),
    .ZN(_14766_));
 OAI211_X1 _24472_ (.A(_14762_),
    .B(_14765_),
    .C1(_14766_),
    .C2(_14672_),
    .ZN(_14767_));
 AND2_X1 _24473_ (.A1(_14700_),
    .A2(_14707_),
    .ZN(_14768_));
 NAND2_X1 _24474_ (.A1(_14768_),
    .A2(_14691_),
    .ZN(_14769_));
 CLKBUF_X2 _24475_ (.A(_14677_),
    .Z(_14770_));
 NAND3_X1 _24476_ (.A1(_14691_),
    .A2(_14708_),
    .A3(_14770_),
    .ZN(_14771_));
 NAND2_X1 _24477_ (.A1(_14769_),
    .A2(_14771_),
    .ZN(_14772_));
 CLKBUF_X2 _24478_ (.A(_14718_),
    .Z(_14773_));
 AND3_X1 _24479_ (.A1(_14691_),
    .A2(_14773_),
    .A3(_14732_),
    .ZN(_14774_));
 NOR4_X1 _24480_ (.A1(_14758_),
    .A2(_14767_),
    .A3(_14772_),
    .A4(_14774_),
    .ZN(_14775_));
 AND2_X1 _24481_ (.A1(_14735_),
    .A2(_14677_),
    .ZN(_14776_));
 BUF_X2 _24482_ (.A(_14776_),
    .Z(_14777_));
 AND2_X1 _24483_ (.A1(_14688_),
    .A2(_14694_),
    .ZN(_14778_));
 BUF_X2 _24484_ (.A(_14778_),
    .Z(_14779_));
 AND2_X1 _24485_ (.A1(_14777_),
    .A2(_14779_),
    .ZN(_14780_));
 BUF_X2 _24486_ (.A(_14698_),
    .Z(_14781_));
 AND2_X2 _24487_ (.A1(_14731_),
    .A2(_14677_),
    .ZN(_14782_));
 BUF_X2 _24488_ (.A(_14734_),
    .Z(_14783_));
 AND2_X1 _24489_ (.A1(_14745_),
    .A2(_14695_),
    .ZN(_14784_));
 AOI221_X4 _24490_ (.A(_14780_),
    .B1(_14781_),
    .B2(_14782_),
    .C1(_14783_),
    .C2(_14784_),
    .ZN(_14785_));
 NAND4_X1 _24491_ (.A1(_14722_),
    .A2(_14746_),
    .A3(_14775_),
    .A4(_14785_),
    .ZN(_14786_));
 AND2_X2 _24492_ (.A1(_14749_),
    .A2(_14694_),
    .ZN(_14787_));
 BUF_X2 _24493_ (.A(_14787_),
    .Z(_14788_));
 AND2_X1 _24494_ (.A1(_14712_),
    .A2(_14677_),
    .ZN(_14789_));
 INV_X1 _24495_ (.A(_14789_),
    .ZN(_14790_));
 AND2_X1 _24496_ (.A1(_14707_),
    .A2(_14677_),
    .ZN(_14791_));
 INV_X1 _24497_ (.A(_14791_),
    .ZN(_14792_));
 NAND2_X1 _24498_ (.A1(_14790_),
    .A2(_14792_),
    .ZN(_14793_));
 AND2_X1 _24499_ (.A1(_14709_),
    .A2(_17067_),
    .ZN(_14794_));
 OAI21_X1 _24500_ (.A(_14788_),
    .B1(_14793_),
    .B2(_14794_),
    .ZN(_14795_));
 CLKBUF_X2 _24501_ (.A(_14791_),
    .Z(_14796_));
 AND2_X1 _24502_ (.A1(_14705_),
    .A2(_14796_),
    .ZN(_14797_));
 INV_X1 _24503_ (.A(_14797_),
    .ZN(_14798_));
 NAND2_X1 _24504_ (.A1(_14795_),
    .A2(_14798_),
    .ZN(_14799_));
 AND2_X1 _24505_ (.A1(_14731_),
    .A2(_14709_),
    .ZN(_14800_));
 CLKBUF_X2 _24506_ (.A(_14800_),
    .Z(_14801_));
 OAI21_X1 _24507_ (.A(_14675_),
    .B1(_14801_),
    .B2(_14687_),
    .ZN(_14802_));
 BUF_X2 _24508_ (.A(_14662_),
    .Z(_14803_));
 NAND4_X1 _24509_ (.A1(_14803_),
    .A2(_04121_),
    .A3(_14701_),
    .A4(_14673_),
    .ZN(_14804_));
 INV_X1 _24510_ (.A(_14681_),
    .ZN(_14805_));
 INV_X1 _24511_ (.A(_14787_),
    .ZN(_14806_));
 OAI211_X1 _24512_ (.A(_14802_),
    .B(_14804_),
    .C1(_14805_),
    .C2(_14806_),
    .ZN(_14807_));
 INV_X1 _24513_ (.A(_14710_),
    .ZN(_14808_));
 AND3_X1 _24514_ (.A1(_14808_),
    .A2(_14781_),
    .A3(_14739_),
    .ZN(_14809_));
 INV_X1 _24515_ (.A(_14779_),
    .ZN(_14810_));
 INV_X1 _24516_ (.A(_14701_),
    .ZN(_14811_));
 INV_X1 _24517_ (.A(_14763_),
    .ZN(_14812_));
 AOI21_X1 _24518_ (.A(_14810_),
    .B1(_14811_),
    .B2(_14812_),
    .ZN(_14813_));
 NOR4_X1 _24519_ (.A1(_14799_),
    .A2(_14807_),
    .A3(_14809_),
    .A4(_14813_),
    .ZN(_14814_));
 AND2_X1 _24520_ (.A1(_14723_),
    .A2(_14688_),
    .ZN(_14815_));
 CLKBUF_X2 _24521_ (.A(_14815_),
    .Z(_14816_));
 AND2_X1 _24522_ (.A1(_14816_),
    .A2(_14747_),
    .ZN(_14817_));
 INV_X1 _24523_ (.A(_14817_),
    .ZN(_14818_));
 NOR2_X1 _24524_ (.A1(_14726_),
    .A2(_14735_),
    .ZN(_14819_));
 NAND2_X1 _24525_ (.A1(_14816_),
    .A2(_14819_),
    .ZN(_14820_));
 BUF_X2 _24526_ (.A(_14683_),
    .Z(_14821_));
 BUF_X2 _24527_ (.A(_14789_),
    .Z(_14822_));
 NAND2_X1 _24528_ (.A1(_14821_),
    .A2(_14822_),
    .ZN(_14823_));
 NAND3_X1 _24529_ (.A1(_14821_),
    .A2(_14783_),
    .A3(_14745_),
    .ZN(_14824_));
 AND4_X1 _24530_ (.A1(_14818_),
    .A2(_14820_),
    .A3(_14823_),
    .A4(_14824_),
    .ZN(_14825_));
 AND2_X1 _24531_ (.A1(_14749_),
    .A2(_14723_),
    .ZN(_14826_));
 AND2_X1 _24532_ (.A1(_14826_),
    .A2(_14755_),
    .ZN(_14827_));
 NAND2_X1 _24533_ (.A1(_14684_),
    .A2(_14777_),
    .ZN(_14828_));
 NAND2_X1 _24534_ (.A1(_14717_),
    .A2(_14796_),
    .ZN(_14829_));
 NAND2_X1 _24535_ (.A1(_14828_),
    .A2(_14829_),
    .ZN(_14830_));
 AND2_X1 _24536_ (.A1(_14723_),
    .A2(_14673_),
    .ZN(_14831_));
 BUF_X2 _24537_ (.A(_14831_),
    .Z(_14832_));
 AOI211_X1 _24538_ (.A(_14827_),
    .B(_14830_),
    .C1(_14808_),
    .C2(_14832_),
    .ZN(_14833_));
 AND2_X1 _24539_ (.A1(_14755_),
    .A2(_14779_),
    .ZN(_14834_));
 AND2_X1 _24540_ (.A1(_14781_),
    .A2(_14759_),
    .ZN(_14835_));
 AND2_X1 _24541_ (.A1(_14782_),
    .A2(_14703_),
    .ZN(_14836_));
 CLKBUF_X2 _24542_ (.A(_14709_),
    .Z(_14837_));
 AND3_X1 _24543_ (.A1(_14778_),
    .A2(_14732_),
    .A3(_14837_),
    .ZN(_14838_));
 NOR4_X1 _24544_ (.A1(_14834_),
    .A2(_14835_),
    .A3(_14836_),
    .A4(_14838_),
    .ZN(_14839_));
 AND4_X1 _24545_ (.A1(_14814_),
    .A2(_14825_),
    .A3(_14833_),
    .A4(_14839_),
    .ZN(_14840_));
 AND2_X1 _24546_ (.A1(_14750_),
    .A2(_14727_),
    .ZN(_14841_));
 INV_X1 _24547_ (.A(_14841_),
    .ZN(_14842_));
 AND2_X1 _24548_ (.A1(_14708_),
    .A2(_14700_),
    .ZN(_14843_));
 NAND2_X1 _24549_ (.A1(_14843_),
    .A2(_14751_),
    .ZN(_14844_));
 NAND2_X1 _24550_ (.A1(_14842_),
    .A2(_14844_),
    .ZN(_14845_));
 NAND2_X1 _24551_ (.A1(_14821_),
    .A2(_14733_),
    .ZN(_14846_));
 INV_X1 _24552_ (.A(_14732_),
    .ZN(_14847_));
 NAND3_X1 _24553_ (.A1(_14831_),
    .A2(_14718_),
    .A3(_14847_),
    .ZN(_14848_));
 NAND3_X1 _24554_ (.A1(_14753_),
    .A2(_14665_),
    .A3(_14803_),
    .ZN(_14849_));
 BUF_X2 _24555_ (.A(_14665_),
    .Z(_14850_));
 BUF_X2 _24556_ (.A(_14700_),
    .Z(_14851_));
 NAND4_X1 _24557_ (.A1(_14803_),
    .A2(_14850_),
    .A3(_14851_),
    .A4(_04132_),
    .ZN(_14852_));
 NAND4_X1 _24558_ (.A1(_14846_),
    .A2(_14848_),
    .A3(_14849_),
    .A4(_14852_),
    .ZN(_14853_));
 AND2_X1 _24559_ (.A1(_14735_),
    .A2(_14709_),
    .ZN(_14854_));
 OAI21_X1 _24560_ (.A(_14716_),
    .B1(_14801_),
    .B2(_14854_),
    .ZN(_14855_));
 AND2_X1 _24561_ (.A1(_14700_),
    .A2(_14712_),
    .ZN(_14856_));
 CLKBUF_X2 _24562_ (.A(_14856_),
    .Z(_14857_));
 CLKBUF_X2 _24563_ (.A(_14688_),
    .Z(_14858_));
 NAND3_X1 _24564_ (.A1(_14857_),
    .A2(_14858_),
    .A3(_14803_),
    .ZN(_14859_));
 NAND2_X1 _24565_ (.A1(_14855_),
    .A2(_14859_),
    .ZN(_14860_));
 NAND2_X1 _24566_ (.A1(_14847_),
    .A2(_14770_),
    .ZN(_14861_));
 NOR2_X1 _24567_ (.A1(_14667_),
    .A2(_14861_),
    .ZN(_14862_));
 NOR4_X1 _24568_ (.A1(_14845_),
    .A2(_14853_),
    .A3(_14860_),
    .A4(_14862_),
    .ZN(_14863_));
 NAND3_X1 _24569_ (.A1(_14787_),
    .A2(_14736_),
    .A3(_14701_),
    .ZN(_14864_));
 CLKBUF_X2 _24570_ (.A(_14826_),
    .Z(_14865_));
 OAI21_X1 _24571_ (.A(_14865_),
    .B1(_14761_),
    .B2(_14687_),
    .ZN(_14866_));
 CLKBUF_X2 _24572_ (.A(_14723_),
    .Z(_14867_));
 NAND4_X1 _24573_ (.A1(_14847_),
    .A2(_14773_),
    .A3(_14858_),
    .A4(_14867_),
    .ZN(_14868_));
 NAND2_X1 _24574_ (.A1(_14865_),
    .A2(_14753_),
    .ZN(_14869_));
 AND4_X1 _24575_ (.A1(_14864_),
    .A2(_14866_),
    .A3(_14868_),
    .A4(_14869_),
    .ZN(_14870_));
 OAI21_X1 _24576_ (.A(_14751_),
    .B1(_14741_),
    .B2(_14745_),
    .ZN(_14871_));
 AND2_X1 _24577_ (.A1(_14770_),
    .A2(_14734_),
    .ZN(_14872_));
 OAI21_X1 _24578_ (.A(_14832_),
    .B1(_14702_),
    .B2(_14872_),
    .ZN(_14873_));
 AND2_X1 _24579_ (.A1(_14871_),
    .A2(_14873_),
    .ZN(_14874_));
 NAND4_X1 _24580_ (.A1(_14840_),
    .A2(_14863_),
    .A3(_14870_),
    .A4(_14874_),
    .ZN(_14875_));
 NOR2_X1 _24581_ (.A1(_14786_),
    .A2(_14875_),
    .ZN(_14876_));
 XOR2_X1 _24582_ (.A(_14876_),
    .B(_00997_),
    .Z(_14877_));
 MUX2_X1 _24583_ (.A(_01207_),
    .B(_14877_),
    .S(_14285_),
    .Z(_01088_));
 INV_X1 _24584_ (.A(_14720_),
    .ZN(_14878_));
 AOI21_X1 _24585_ (.A(_14676_),
    .B1(_14878_),
    .B2(_14740_),
    .ZN(_14879_));
 INV_X1 _24586_ (.A(_14709_),
    .ZN(_14880_));
 AOI211_X1 _24587_ (.A(_14880_),
    .B(_14676_),
    .C1(_14847_),
    .C2(_14736_),
    .ZN(_14881_));
 AOI211_X1 _24588_ (.A(_14879_),
    .B(_14881_),
    .C1(_14851_),
    .C2(_14675_),
    .ZN(_14882_));
 CLKBUF_X2 _24589_ (.A(_14666_),
    .Z(_14883_));
 AND2_X2 _24590_ (.A1(_14700_),
    .A2(_09451_),
    .ZN(_14884_));
 AND2_X1 _24591_ (.A1(_14883_),
    .A2(_14884_),
    .ZN(_14885_));
 INV_X1 _24592_ (.A(_14885_),
    .ZN(_14886_));
 AND2_X1 _24593_ (.A1(_14669_),
    .A2(_14712_),
    .ZN(_14887_));
 CLKBUF_X2 _24594_ (.A(_14887_),
    .Z(_14888_));
 OAI211_X1 _24595_ (.A(_14850_),
    .B(_14803_),
    .C1(_14888_),
    .C2(_14796_),
    .ZN(_14889_));
 OAI211_X1 _24596_ (.A(_14850_),
    .B(_14803_),
    .C1(_14753_),
    .C2(_14748_),
    .ZN(_14890_));
 AND2_X1 _24597_ (.A1(_14731_),
    .A2(_14700_),
    .ZN(_14891_));
 CLKBUF_X2 _24598_ (.A(_14891_),
    .Z(_14892_));
 NAND3_X1 _24599_ (.A1(_14892_),
    .A2(_14850_),
    .A3(_14803_),
    .ZN(_14893_));
 AND4_X1 _24600_ (.A1(_14886_),
    .A2(_14889_),
    .A3(_14890_),
    .A4(_14893_),
    .ZN(_14894_));
 NAND2_X1 _24601_ (.A1(_14708_),
    .A2(_14770_),
    .ZN(_14895_));
 INV_X1 _24602_ (.A(_14895_),
    .ZN(_14896_));
 AND2_X1 _24603_ (.A1(_14896_),
    .A2(_14684_),
    .ZN(_14897_));
 NAND2_X1 _24604_ (.A1(_14684_),
    .A2(_14801_),
    .ZN(_14898_));
 INV_X1 _24605_ (.A(_14714_),
    .ZN(_14899_));
 OAI21_X1 _24606_ (.A(_14898_),
    .B1(_14757_),
    .B2(_14899_),
    .ZN(_14900_));
 AND2_X1 _24607_ (.A1(_14718_),
    .A2(_14734_),
    .ZN(_14901_));
 AOI211_X1 _24608_ (.A(_14897_),
    .B(_14900_),
    .C1(_14901_),
    .C2(_14821_),
    .ZN(_14902_));
 AND2_X1 _24609_ (.A1(_14808_),
    .A2(_14716_),
    .ZN(_14903_));
 INV_X1 _24610_ (.A(_14716_),
    .ZN(_14904_));
 AOI21_X1 _24611_ (.A(_14904_),
    .B1(_14756_),
    .B2(_14878_),
    .ZN(_14905_));
 AND2_X1 _24612_ (.A1(_14843_),
    .A2(_14739_),
    .ZN(_14906_));
 AOI211_X1 _24613_ (.A(_14903_),
    .B(_14905_),
    .C1(_14717_),
    .C2(_14906_),
    .ZN(_14907_));
 AND4_X1 _24614_ (.A1(_14882_),
    .A2(_14894_),
    .A3(_14902_),
    .A4(_14907_),
    .ZN(_14908_));
 AND2_X1 _24615_ (.A1(_14698_),
    .A2(_14747_),
    .ZN(_14909_));
 AND2_X1 _24616_ (.A1(_14698_),
    .A2(_14892_),
    .ZN(_14910_));
 AOI211_X1 _24617_ (.A(_14909_),
    .B(_14910_),
    .C1(_14781_),
    .C2(_14753_),
    .ZN(_14911_));
 OAI21_X1 _24618_ (.A(_14781_),
    .B1(_14760_),
    .B2(_14671_),
    .ZN(_14912_));
 INV_X1 _24619_ (.A(_14698_),
    .ZN(_14913_));
 OAI211_X1 _24620_ (.A(_14911_),
    .B(_14912_),
    .C1(_14913_),
    .C2(_14878_),
    .ZN(_14914_));
 OAI21_X1 _24621_ (.A(_14695_),
    .B1(_14789_),
    .B2(_14791_),
    .ZN(_14915_));
 INV_X1 _24622_ (.A(_14719_),
    .ZN(_14916_));
 INV_X1 _24623_ (.A(_14695_),
    .ZN(_14917_));
 OAI21_X1 _24624_ (.A(_14915_),
    .B1(_14916_),
    .B2(_14917_),
    .ZN(_14918_));
 AND2_X1 _24625_ (.A1(_14857_),
    .A2(_14695_),
    .ZN(_14919_));
 AND2_X1 _24626_ (.A1(_14747_),
    .A2(_14695_),
    .ZN(_14920_));
 OR4_X1 _24627_ (.A1(_14784_),
    .A2(_14918_),
    .A3(_14919_),
    .A4(_14920_),
    .ZN(_14921_));
 AND2_X1 _24628_ (.A1(_14788_),
    .A2(_14884_),
    .ZN(_14922_));
 INV_X1 _24629_ (.A(_14922_),
    .ZN(_14923_));
 AND2_X2 _24630_ (.A1(_14718_),
    .A2(_14731_),
    .ZN(_14924_));
 AND2_X1 _24631_ (.A1(_14924_),
    .A2(_14787_),
    .ZN(_14925_));
 INV_X1 _24632_ (.A(_14925_),
    .ZN(_14926_));
 NAND2_X1 _24633_ (.A1(_14892_),
    .A2(_14788_),
    .ZN(_14927_));
 OAI21_X1 _24634_ (.A(_14787_),
    .B1(_14753_),
    .B2(_14747_),
    .ZN(_14928_));
 NAND4_X1 _24635_ (.A1(_14923_),
    .A2(_14926_),
    .A3(_14927_),
    .A4(_14928_),
    .ZN(_14929_));
 AND2_X1 _24636_ (.A1(_14681_),
    .A2(_14778_),
    .ZN(_14930_));
 INV_X1 _24637_ (.A(_14930_),
    .ZN(_14931_));
 NAND2_X1 _24638_ (.A1(_14779_),
    .A2(_14745_),
    .ZN(_14932_));
 NAND2_X1 _24639_ (.A1(_14857_),
    .A2(_14779_),
    .ZN(_14933_));
 NAND2_X1 _24640_ (.A1(_14924_),
    .A2(_14779_),
    .ZN(_14934_));
 NAND4_X1 _24641_ (.A1(_14931_),
    .A2(_14932_),
    .A3(_14933_),
    .A4(_14934_),
    .ZN(_14935_));
 NOR4_X1 _24642_ (.A1(_14914_),
    .A2(_14921_),
    .A3(_14929_),
    .A4(_14935_),
    .ZN(_14936_));
 AND2_X1 _24643_ (.A1(_14714_),
    .A2(_14705_),
    .ZN(_14937_));
 AOI21_X1 _24644_ (.A(_14766_),
    .B1(_14740_),
    .B2(_14812_),
    .ZN(_14938_));
 AOI211_X1 _24645_ (.A(_14937_),
    .B(_14938_),
    .C1(_14837_),
    .C2(_14706_),
    .ZN(_14939_));
 INV_X1 _24646_ (.A(_14901_),
    .ZN(_14940_));
 AOI21_X1 _24647_ (.A(_14730_),
    .B1(_14679_),
    .B2(_14940_),
    .ZN(_14941_));
 CLKBUF_X2 _24648_ (.A(_14729_),
    .Z(_14942_));
 AND2_X1 _24649_ (.A1(_14942_),
    .A2(_14801_),
    .ZN(_14943_));
 AND2_X1 _24650_ (.A1(_14729_),
    .A2(_14714_),
    .ZN(_14944_));
 NOR3_X1 _24651_ (.A1(_14941_),
    .A2(_14943_),
    .A3(_14944_),
    .ZN(_14945_));
 INV_X1 _24652_ (.A(_14750_),
    .ZN(_14946_));
 NOR2_X1 _24653_ (.A1(_14946_),
    .A2(_14740_),
    .ZN(_14947_));
 AOI21_X1 _24654_ (.A(_14947_),
    .B1(_14751_),
    .B2(_14819_),
    .ZN(_14948_));
 NAND2_X1 _24655_ (.A1(_14691_),
    .A2(_14687_),
    .ZN(_14949_));
 OAI21_X1 _24656_ (.A(_14690_),
    .B1(_14896_),
    .B2(_14719_),
    .ZN(_14950_));
 NAND2_X1 _24657_ (.A1(_14801_),
    .A2(_14690_),
    .ZN(_14951_));
 OAI211_X1 _24658_ (.A(_14690_),
    .B(_14701_),
    .C1(_04121_),
    .C2(_09452_),
    .ZN(_14952_));
 AND4_X1 _24659_ (.A1(_14949_),
    .A2(_14950_),
    .A3(_14951_),
    .A4(_14952_),
    .ZN(_14953_));
 AND4_X1 _24660_ (.A1(_14939_),
    .A2(_14945_),
    .A3(_14948_),
    .A4(_14953_),
    .ZN(_14954_));
 OAI211_X1 _24661_ (.A(_14816_),
    .B(_14837_),
    .C1(_14732_),
    .C2(_14735_),
    .ZN(_14955_));
 BUF_X2 _24662_ (.A(_14816_),
    .Z(_14956_));
 OAI21_X1 _24663_ (.A(_14956_),
    .B1(_14924_),
    .B2(_14872_),
    .ZN(_14957_));
 NAND4_X1 _24664_ (.A1(_14851_),
    .A2(_14867_),
    .A3(_04121_),
    .A4(_14858_),
    .ZN(_14958_));
 AND3_X1 _24665_ (.A1(_14955_),
    .A2(_14957_),
    .A3(_14958_),
    .ZN(_14959_));
 AND2_X1 _24666_ (.A1(_14725_),
    .A2(_14837_),
    .ZN(_14960_));
 NAND3_X1 _24667_ (.A1(_14782_),
    .A2(_14665_),
    .A3(_14867_),
    .ZN(_14961_));
 INV_X2 _24668_ (.A(_14724_),
    .ZN(_14962_));
 OAI21_X1 _24669_ (.A(_14961_),
    .B1(_14962_),
    .B2(_14805_),
    .ZN(_14963_));
 AOI211_X1 _24670_ (.A(_14960_),
    .B(_14963_),
    .C1(_14884_),
    .C2(_14725_),
    .ZN(_14964_));
 AND3_X1 _24671_ (.A1(_14843_),
    .A2(_14739_),
    .A3(_14831_),
    .ZN(_14965_));
 NAND4_X1 _24672_ (.A1(_14732_),
    .A2(_14867_),
    .A3(_14673_),
    .A4(_14770_),
    .ZN(_14966_));
 NAND2_X1 _24673_ (.A1(_14848_),
    .A2(_14966_),
    .ZN(_14967_));
 AOI211_X1 _24674_ (.A(_14965_),
    .B(_14967_),
    .C1(_14832_),
    .C2(_14753_),
    .ZN(_14968_));
 AND2_X1 _24675_ (.A1(_14865_),
    .A2(_14763_),
    .ZN(_14969_));
 AND2_X1 _24676_ (.A1(_14759_),
    .A2(_14865_),
    .ZN(_14970_));
 AND2_X1 _24677_ (.A1(_14733_),
    .A2(_14826_),
    .ZN(_14971_));
 AND2_X1 _24678_ (.A1(_14865_),
    .A2(_14777_),
    .ZN(_14972_));
 NOR4_X1 _24679_ (.A1(_14969_),
    .A2(_14970_),
    .A3(_14971_),
    .A4(_14972_),
    .ZN(_14973_));
 AND4_X1 _24680_ (.A1(_14959_),
    .A2(_14964_),
    .A3(_14968_),
    .A4(_14973_),
    .ZN(_14974_));
 NAND4_X1 _24681_ (.A1(_14908_),
    .A2(_14936_),
    .A3(_14954_),
    .A4(_14974_),
    .ZN(_14975_));
 NOR2_X1 _24682_ (.A1(_14975_),
    .A2(_14797_),
    .ZN(_14976_));
 INV_X1 _24683_ (.A(_00998_),
    .ZN(_14977_));
 XNOR2_X1 _24684_ (.A(_14976_),
    .B(_14977_),
    .ZN(_14978_));
 MUX2_X1 _24685_ (.A(_01208_),
    .B(_14978_),
    .S(_14285_),
    .Z(_01089_));
 OAI21_X1 _24686_ (.A(_14821_),
    .B1(_14737_),
    .B2(_14713_),
    .ZN(_14979_));
 AND2_X1 _24687_ (.A1(_14683_),
    .A2(_14888_),
    .ZN(_14980_));
 AND2_X1 _24688_ (.A1(_14683_),
    .A2(_14678_),
    .ZN(_14981_));
 AOI221_X4 _24689_ (.A(_14980_),
    .B1(_14759_),
    .B2(_14684_),
    .C1(_04121_),
    .C2(_14981_),
    .ZN(_14982_));
 OAI21_X1 _24690_ (.A(_14717_),
    .B1(_14719_),
    .B2(_14822_),
    .ZN(_14983_));
 BUF_X2 _24691_ (.A(_14854_),
    .Z(_14984_));
 OAI21_X1 _24692_ (.A(_14717_),
    .B1(_14984_),
    .B2(_14884_),
    .ZN(_14985_));
 AND4_X1 _24693_ (.A1(_14979_),
    .A2(_14982_),
    .A3(_14983_),
    .A4(_14985_),
    .ZN(_14986_));
 NAND2_X1 _24694_ (.A1(_14847_),
    .A2(_14709_),
    .ZN(_14987_));
 INV_X1 _24695_ (.A(_14987_),
    .ZN(_14988_));
 NAND2_X1 _24696_ (.A1(_14988_),
    .A2(_14706_),
    .ZN(_14989_));
 NAND3_X1 _24697_ (.A1(_14706_),
    .A2(_14732_),
    .A3(_14851_),
    .ZN(_14990_));
 AND2_X1 _24698_ (.A1(_14989_),
    .A2(_14990_),
    .ZN(_14991_));
 AND2_X1 _24699_ (.A1(_14671_),
    .A2(_14705_),
    .ZN(_14992_));
 NAND2_X1 _24700_ (.A1(_14896_),
    .A2(_14705_),
    .ZN(_14993_));
 INV_X1 _24701_ (.A(_14993_),
    .ZN(_14994_));
 AOI21_X1 _24702_ (.A(_14992_),
    .B1(_14994_),
    .B2(_14739_),
    .ZN(_14995_));
 OAI211_X1 _24703_ (.A(_14942_),
    .B(_14851_),
    .C1(_04121_),
    .C2(_09452_),
    .ZN(_14996_));
 NAND3_X1 _24704_ (.A1(_14687_),
    .A2(_14850_),
    .A3(_14764_),
    .ZN(_14997_));
 AND2_X1 _24705_ (.A1(_14996_),
    .A2(_14997_),
    .ZN(_14998_));
 OAI21_X1 _24706_ (.A(_14942_),
    .B1(_14924_),
    .B2(_14822_),
    .ZN(_14999_));
 AND4_X1 _24707_ (.A1(_14991_),
    .A2(_14995_),
    .A3(_14998_),
    .A4(_14999_),
    .ZN(_15000_));
 INV_X1 _24708_ (.A(_14690_),
    .ZN(_15001_));
 AOI21_X1 _24709_ (.A(_15001_),
    .B1(_14742_),
    .B2(_14679_),
    .ZN(_15002_));
 OAI21_X1 _24710_ (.A(_14751_),
    .B1(_14777_),
    .B2(_14796_),
    .ZN(_15003_));
 NAND2_X1 _24711_ (.A1(_14751_),
    .A2(_14681_),
    .ZN(_15004_));
 NAND3_X1 _24712_ (.A1(_14822_),
    .A2(_14749_),
    .A3(_14764_),
    .ZN(_15005_));
 NAND2_X1 _24713_ (.A1(_14751_),
    .A2(_14671_),
    .ZN(_15006_));
 NAND4_X1 _24714_ (.A1(_15003_),
    .A2(_15004_),
    .A3(_15005_),
    .A4(_15006_),
    .ZN(_15007_));
 NAND4_X1 _24715_ (.A1(_14732_),
    .A2(_14851_),
    .A3(_14749_),
    .A4(_14764_),
    .ZN(_15008_));
 NAND4_X1 _24716_ (.A1(_14749_),
    .A2(_14837_),
    .A3(_14712_),
    .A4(_14764_),
    .ZN(_15009_));
 INV_X1 _24717_ (.A(_14884_),
    .ZN(_15010_));
 OAI211_X1 _24718_ (.A(_15008_),
    .B(_15009_),
    .C1(_15010_),
    .C2(_14946_),
    .ZN(_15011_));
 INV_X1 _24719_ (.A(_14768_),
    .ZN(_15012_));
 INV_X1 _24720_ (.A(_14794_),
    .ZN(_15013_));
 AOI21_X1 _24721_ (.A(_15001_),
    .B1(_15012_),
    .B2(_15013_),
    .ZN(_15014_));
 NOR4_X1 _24722_ (.A1(_15002_),
    .A2(_15007_),
    .A3(_15011_),
    .A4(_15014_),
    .ZN(_15015_));
 OAI21_X1 _24723_ (.A(_14675_),
    .B1(_14760_),
    .B2(_14782_),
    .ZN(_15016_));
 OAI21_X1 _24724_ (.A(_14883_),
    .B1(_14760_),
    .B2(_14822_),
    .ZN(_15017_));
 OAI21_X1 _24725_ (.A(_14883_),
    .B1(_14892_),
    .B2(_14794_),
    .ZN(_15018_));
 OAI21_X1 _24726_ (.A(_14675_),
    .B1(_14892_),
    .B2(_14745_),
    .ZN(_15019_));
 AND4_X1 _24727_ (.A1(_15016_),
    .A2(_15017_),
    .A3(_15018_),
    .A4(_15019_),
    .ZN(_15020_));
 NAND4_X1 _24728_ (.A1(_14986_),
    .A2(_15000_),
    .A3(_15015_),
    .A4(_15020_),
    .ZN(_15021_));
 AOI211_X1 _24729_ (.A(_14811_),
    .B(_14917_),
    .C1(_14783_),
    .C2(_09452_),
    .ZN(_15022_));
 AND2_X1 _24730_ (.A1(_14984_),
    .A2(_14703_),
    .ZN(_15023_));
 OR2_X1 _24731_ (.A1(_15022_),
    .A2(_15023_),
    .ZN(_15024_));
 OAI21_X1 _24732_ (.A(_14781_),
    .B1(_14892_),
    .B2(_14761_),
    .ZN(_15025_));
 OAI21_X1 _24733_ (.A(_14781_),
    .B1(_14777_),
    .B2(_14763_),
    .ZN(_15026_));
 OAI211_X1 _24734_ (.A(_14694_),
    .B(_14850_),
    .C1(_14745_),
    .C2(_14748_),
    .ZN(_15027_));
 NAND2_X1 _24735_ (.A1(_14781_),
    .A2(_14671_),
    .ZN(_15028_));
 NAND4_X1 _24736_ (.A1(_15025_),
    .A2(_15026_),
    .A3(_15027_),
    .A4(_15028_),
    .ZN(_15029_));
 AND3_X1 _24737_ (.A1(_14718_),
    .A2(_14694_),
    .A3(_14673_),
    .ZN(_15030_));
 INV_X1 _24738_ (.A(_14782_),
    .ZN(_15031_));
 AOI21_X1 _24739_ (.A(_14917_),
    .B1(_15031_),
    .B2(_14790_),
    .ZN(_15032_));
 NOR4_X1 _24740_ (.A1(_15024_),
    .A2(_15029_),
    .A3(_15030_),
    .A4(_15032_),
    .ZN(_15033_));
 OAI21_X1 _24741_ (.A(_14725_),
    .B1(_14857_),
    .B2(_14884_),
    .ZN(_15034_));
 NAND2_X1 _24742_ (.A1(_14725_),
    .A2(_14763_),
    .ZN(_15035_));
 INV_X1 _24743_ (.A(_14687_),
    .ZN(_15036_));
 OAI211_X1 _24744_ (.A(_15034_),
    .B(_15035_),
    .C1(_15036_),
    .C2(_14962_),
    .ZN(_15037_));
 INV_X1 _24745_ (.A(_14832_),
    .ZN(_15038_));
 NOR2_X1 _24746_ (.A1(_15038_),
    .A2(_14861_),
    .ZN(_15039_));
 NAND2_X1 _24747_ (.A1(_14832_),
    .A2(_14687_),
    .ZN(_15040_));
 OAI21_X1 _24748_ (.A(_15040_),
    .B1(_15038_),
    .B2(_14811_),
    .ZN(_15041_));
 AND2_X1 _24749_ (.A1(_14832_),
    .A2(_14773_),
    .ZN(_15042_));
 NOR4_X1 _24750_ (.A1(_15037_),
    .A2(_15039_),
    .A3(_15041_),
    .A4(_15042_),
    .ZN(_15043_));
 OAI21_X1 _24751_ (.A(_14865_),
    .B1(_14713_),
    .B2(_14892_),
    .ZN(_15044_));
 NAND2_X1 _24752_ (.A1(_14760_),
    .A2(_14865_),
    .ZN(_15045_));
 NAND2_X1 _24753_ (.A1(_14865_),
    .A2(_14671_),
    .ZN(_15046_));
 AND3_X1 _24754_ (.A1(_15044_),
    .A2(_15045_),
    .A3(_15046_),
    .ZN(_15047_));
 OAI211_X1 _24755_ (.A(_14956_),
    .B(_14773_),
    .C1(_14783_),
    .C2(_09452_),
    .ZN(_15048_));
 OAI211_X1 _24756_ (.A(_14816_),
    .B(_14701_),
    .C1(_14783_),
    .C2(_09452_),
    .ZN(_15049_));
 OAI21_X1 _24757_ (.A(_14816_),
    .B1(_14801_),
    .B2(_14748_),
    .ZN(_15050_));
 AND2_X1 _24758_ (.A1(_15049_),
    .A2(_15050_),
    .ZN(_15051_));
 AND4_X1 _24759_ (.A1(_14820_),
    .A2(_15047_),
    .A3(_15048_),
    .A4(_15051_),
    .ZN(_15052_));
 NAND2_X1 _24760_ (.A1(_14788_),
    .A2(_14671_),
    .ZN(_15053_));
 AND4_X1 _24761_ (.A1(_14778_),
    .A2(_14847_),
    .A3(_14736_),
    .A4(_14770_),
    .ZN(_15054_));
 AND2_X1 _24762_ (.A1(_14714_),
    .A2(_14778_),
    .ZN(_15055_));
 AND4_X1 _24763_ (.A1(_04121_),
    .A2(_14858_),
    .A3(_14694_),
    .A4(_14709_),
    .ZN(_15056_));
 NOR4_X1 _24764_ (.A1(_14930_),
    .A2(_15054_),
    .A3(_15055_),
    .A4(_15056_),
    .ZN(_15057_));
 AND2_X1 _24765_ (.A1(_14787_),
    .A2(_14794_),
    .ZN(_15058_));
 AND2_X1 _24766_ (.A1(_14787_),
    .A2(_14747_),
    .ZN(_15059_));
 NOR2_X1 _24767_ (.A1(_15058_),
    .A2(_15059_),
    .ZN(_15060_));
 NAND3_X1 _24768_ (.A1(_14843_),
    .A2(_14788_),
    .A3(_14739_),
    .ZN(_15061_));
 AND4_X1 _24769_ (.A1(_15053_),
    .A2(_15057_),
    .A3(_15060_),
    .A4(_15061_),
    .ZN(_15062_));
 NAND4_X1 _24770_ (.A1(_15033_),
    .A2(_15043_),
    .A3(_15052_),
    .A4(_15062_),
    .ZN(_15063_));
 NOR2_X1 _24771_ (.A1(_15021_),
    .A2(_15063_),
    .ZN(_15064_));
 XOR2_X1 _24772_ (.A(_15064_),
    .B(_00999_),
    .Z(_15065_));
 MUX2_X1 _24773_ (.A(_01209_),
    .B(_15065_),
    .S(_14285_),
    .Z(_01059_));
 NAND4_X1 _24774_ (.A1(_14867_),
    .A2(_04132_),
    .A3(_14858_),
    .A4(_14770_),
    .ZN(_15066_));
 AND2_X1 _24775_ (.A1(_14892_),
    .A2(_14826_),
    .ZN(_15067_));
 INV_X1 _24776_ (.A(_15067_),
    .ZN(_15068_));
 NAND2_X1 _24777_ (.A1(_15068_),
    .A2(_14869_),
    .ZN(_15069_));
 AND2_X1 _24778_ (.A1(_14826_),
    .A2(_14888_),
    .ZN(_15070_));
 NOR4_X1 _24779_ (.A1(_15069_),
    .A2(_14827_),
    .A3(_14969_),
    .A4(_15070_),
    .ZN(_15071_));
 OAI211_X1 _24780_ (.A(_14956_),
    .B(_14773_),
    .C1(_14783_),
    .C2(_09041_),
    .ZN(_15072_));
 AND4_X1 _24781_ (.A1(_09041_),
    .A2(_14867_),
    .A3(_14858_),
    .A4(_14837_),
    .ZN(_15073_));
 AND2_X1 _24782_ (.A1(_14984_),
    .A2(_14816_),
    .ZN(_15074_));
 AOI211_X1 _24783_ (.A(_15073_),
    .B(_15074_),
    .C1(_14956_),
    .C2(_14737_),
    .ZN(_15075_));
 AND4_X1 _24784_ (.A1(_15066_),
    .A2(_15071_),
    .A3(_15072_),
    .A4(_15075_),
    .ZN(_15076_));
 OAI21_X1 _24785_ (.A(_14832_),
    .B1(_14713_),
    .B2(_14714_),
    .ZN(_15077_));
 NAND2_X1 _24786_ (.A1(_14755_),
    .A2(_14832_),
    .ZN(_15078_));
 OAI211_X1 _24787_ (.A(_15077_),
    .B(_15078_),
    .C1(_15038_),
    .C2(_14861_),
    .ZN(_15079_));
 AND2_X1 _24788_ (.A1(_14906_),
    .A2(_14725_),
    .ZN(_15080_));
 OAI21_X1 _24789_ (.A(_15035_),
    .B1(_14962_),
    .B2(_14916_),
    .ZN(_15081_));
 NOR4_X1 _24790_ (.A1(_15079_),
    .A2(_15080_),
    .A3(_14960_),
    .A4(_15081_),
    .ZN(_15082_));
 NAND3_X1 _24791_ (.A1(_14703_),
    .A2(_14773_),
    .A3(_14707_),
    .ZN(_15083_));
 INV_X1 _24792_ (.A(_14887_),
    .ZN(_15084_));
 AOI21_X1 _24793_ (.A(_14913_),
    .B1(_14756_),
    .B2(_15084_),
    .ZN(_15085_));
 AND2_X1 _24794_ (.A1(_14697_),
    .A2(_14857_),
    .ZN(_15086_));
 AND2_X1 _24795_ (.A1(_14698_),
    .A2(_14745_),
    .ZN(_15087_));
 AND3_X1 _24796_ (.A1(_14776_),
    .A2(_14694_),
    .A3(_14665_),
    .ZN(_15088_));
 NOR4_X1 _24797_ (.A1(_15085_),
    .A2(_15086_),
    .A3(_15087_),
    .A4(_15088_),
    .ZN(_15089_));
 AND2_X1 _24798_ (.A1(_14884_),
    .A2(_14695_),
    .ZN(_15090_));
 NOR4_X1 _24799_ (.A1(_14919_),
    .A2(_15090_),
    .A3(_14784_),
    .A4(_14696_),
    .ZN(_15091_));
 OAI21_X1 _24800_ (.A(_14703_),
    .B1(_14822_),
    .B2(_14678_),
    .ZN(_15092_));
 AND4_X1 _24801_ (.A1(_15083_),
    .A2(_15089_),
    .A3(_15091_),
    .A4(_15092_),
    .ZN(_15093_));
 AND2_X1 _24802_ (.A1(_14761_),
    .A2(_14778_),
    .ZN(_15094_));
 NOR3_X1 _24803_ (.A1(_15055_),
    .A2(_15094_),
    .A3(_14838_),
    .ZN(_15095_));
 INV_X1 _24804_ (.A(_14834_),
    .ZN(_15096_));
 AND2_X1 _24805_ (.A1(_14888_),
    .A2(_14778_),
    .ZN(_15097_));
 INV_X1 _24806_ (.A(_15097_),
    .ZN(_15098_));
 OAI21_X1 _24807_ (.A(_14779_),
    .B1(_14796_),
    .B2(_14763_),
    .ZN(_15099_));
 NAND4_X1 _24808_ (.A1(_15095_),
    .A2(_15096_),
    .A3(_15098_),
    .A4(_15099_),
    .ZN(_15100_));
 INV_X1 _24809_ (.A(_14777_),
    .ZN(_15101_));
 AOI21_X1 _24810_ (.A(_14806_),
    .B1(_15031_),
    .B2(_15101_),
    .ZN(_15102_));
 INV_X1 _24811_ (.A(_14924_),
    .ZN(_15103_));
 AOI21_X1 _24812_ (.A(_14806_),
    .B1(_14805_),
    .B2(_15103_),
    .ZN(_15104_));
 OAI21_X1 _24813_ (.A(_14788_),
    .B1(_14748_),
    .B2(_14745_),
    .ZN(_15105_));
 NAND2_X1 _24814_ (.A1(_14788_),
    .A2(_14857_),
    .ZN(_15106_));
 OAI211_X1 _24815_ (.A(_15105_),
    .B(_15106_),
    .C1(_14806_),
    .C2(_15010_),
    .ZN(_15107_));
 NOR4_X1 _24816_ (.A1(_15100_),
    .A2(_15102_),
    .A3(_15104_),
    .A4(_15107_),
    .ZN(_15108_));
 NAND4_X1 _24817_ (.A1(_15076_),
    .A2(_15082_),
    .A3(_15093_),
    .A4(_15108_),
    .ZN(_15109_));
 OAI21_X1 _24818_ (.A(_14821_),
    .B1(_14896_),
    .B2(_14760_),
    .ZN(_15110_));
 AND3_X1 _24819_ (.A1(_14854_),
    .A2(_14749_),
    .A3(_14803_),
    .ZN(_15111_));
 AND2_X1 _24820_ (.A1(_14684_),
    .A2(_14702_),
    .ZN(_15112_));
 AOI211_X1 _24821_ (.A(_15111_),
    .B(_15112_),
    .C1(_14745_),
    .C2(_14821_),
    .ZN(_15113_));
 OAI21_X1 _24822_ (.A(_14717_),
    .B1(_14741_),
    .B2(_14822_),
    .ZN(_15114_));
 AND2_X1 _24823_ (.A1(_14701_),
    .A2(_14734_),
    .ZN(_15115_));
 OAI21_X1 _24824_ (.A(_14717_),
    .B1(_14984_),
    .B2(_15115_),
    .ZN(_15116_));
 AND4_X1 _24825_ (.A1(_15110_),
    .A2(_15113_),
    .A3(_15114_),
    .A4(_15116_),
    .ZN(_15117_));
 NAND3_X1 _24826_ (.A1(_14748_),
    .A2(_14850_),
    .A3(_14764_),
    .ZN(_15118_));
 OAI21_X1 _24827_ (.A(_15118_),
    .B1(_14738_),
    .B2(_14730_),
    .ZN(_15119_));
 OAI21_X1 _24828_ (.A(_14942_),
    .B1(_14782_),
    .B2(_14822_),
    .ZN(_15120_));
 NAND4_X1 _24829_ (.A1(_14850_),
    .A2(_14707_),
    .A3(_14764_),
    .A4(_14770_),
    .ZN(_15121_));
 OAI211_X1 _24830_ (.A(_15120_),
    .B(_15121_),
    .C1(_14805_),
    .C2(_14730_),
    .ZN(_15122_));
 AOI21_X1 _24831_ (.A(_14766_),
    .B1(_14742_),
    .B2(_14878_),
    .ZN(_15123_));
 NAND2_X1 _24832_ (.A1(_14801_),
    .A2(_14706_),
    .ZN(_15124_));
 NAND3_X1 _24833_ (.A1(_14706_),
    .A2(_14712_),
    .A3(_14851_),
    .ZN(_15125_));
 NAND2_X1 _24834_ (.A1(_14687_),
    .A2(_14706_),
    .ZN(_15126_));
 OAI211_X1 _24835_ (.A(_15124_),
    .B(_15125_),
    .C1(_04132_),
    .C2(_15126_),
    .ZN(_15127_));
 NOR4_X1 _24836_ (.A1(_15119_),
    .A2(_15122_),
    .A3(_15123_),
    .A4(_15127_),
    .ZN(_15128_));
 NAND2_X1 _24837_ (.A1(_14984_),
    .A2(_14751_),
    .ZN(_15129_));
 OAI21_X1 _24838_ (.A(_14691_),
    .B1(_14755_),
    .B2(_14888_),
    .ZN(_15130_));
 OAI21_X1 _24839_ (.A(_14751_),
    .B1(_14777_),
    .B2(_14719_),
    .ZN(_15131_));
 NAND2_X1 _24840_ (.A1(_14748_),
    .A2(_14691_),
    .ZN(_15132_));
 AND4_X1 _24841_ (.A1(_15129_),
    .A2(_15130_),
    .A3(_15131_),
    .A4(_15132_),
    .ZN(_15133_));
 OAI211_X1 _24842_ (.A(_14675_),
    .B(_14770_),
    .C1(_14783_),
    .C2(_09041_),
    .ZN(_15134_));
 AND2_X1 _24843_ (.A1(_14709_),
    .A2(_14734_),
    .ZN(_15135_));
 OAI21_X1 _24844_ (.A(_14675_),
    .B1(_14761_),
    .B2(_15135_),
    .ZN(_15136_));
 OAI211_X1 _24845_ (.A(_15134_),
    .B(_15136_),
    .C1(_14676_),
    .C2(_14740_),
    .ZN(_15137_));
 OAI211_X1 _24846_ (.A(_14665_),
    .B(_14662_),
    .C1(_14800_),
    .C2(_14752_),
    .ZN(_15138_));
 OAI21_X1 _24847_ (.A(_15138_),
    .B1(_15036_),
    .B2(_14667_),
    .ZN(_15139_));
 AOI21_X1 _24848_ (.A(_14667_),
    .B1(_15010_),
    .B2(_14899_),
    .ZN(_15140_));
 NAND2_X1 _24849_ (.A1(_14883_),
    .A2(_14719_),
    .ZN(_15141_));
 OAI21_X1 _24850_ (.A(_15141_),
    .B1(_14667_),
    .B2(_14790_),
    .ZN(_15142_));
 NOR4_X1 _24851_ (.A1(_15137_),
    .A2(_15139_),
    .A3(_15140_),
    .A4(_15142_),
    .ZN(_15143_));
 NAND4_X1 _24852_ (.A1(_15117_),
    .A2(_15128_),
    .A3(_15133_),
    .A4(_15143_),
    .ZN(_15144_));
 NOR2_X1 _24853_ (.A1(_15109_),
    .A2(_15144_),
    .ZN(_15145_));
 XOR2_X1 _24854_ (.A(_15145_),
    .B(_01000_),
    .Z(_15146_));
 BUF_X2 _24855_ (.A(_03738_),
    .Z(_15147_));
 MUX2_X1 _24856_ (.A(_01210_),
    .B(_15146_),
    .S(_15147_),
    .Z(_01060_));
 XOR2_X1 _24857_ (.A(_17194_),
    .B(_16998_),
    .Z(_15148_));
 XOR2_X2 _24858_ (.A(_11548_),
    .B(_13842_),
    .Z(_15149_));
 XNOR2_X1 _24859_ (.A(_12285_),
    .B(_15149_),
    .ZN(_15150_));
 XNOR2_X1 _24860_ (.A(_12500_),
    .B(_12807_),
    .ZN(_15151_));
 XNOR2_X1 _24861_ (.A(_15150_),
    .B(_15151_),
    .ZN(_15152_));
 INV_X1 _24862_ (.A(_17194_),
    .ZN(_15153_));
 XNOR2_X1 _24863_ (.A(_15152_),
    .B(_15153_),
    .ZN(_15154_));
 BUF_X2 _24864_ (.A(_09039_),
    .Z(_15155_));
 MUX2_X1 _24865_ (.A(_15148_),
    .B(_15154_),
    .S(_15155_),
    .Z(_00685_));
 INV_X1 _24866_ (.A(_14744_),
    .ZN(_15156_));
 AOI211_X1 _24867_ (.A(_04132_),
    .B(_14730_),
    .C1(_15156_),
    .C2(_15036_),
    .ZN(_15157_));
 AND2_X1 _24868_ (.A1(_14942_),
    .A2(_14789_),
    .ZN(_15158_));
 AND2_X1 _24869_ (.A1(_14729_),
    .A2(_14761_),
    .ZN(_15159_));
 AOI21_X1 _24870_ (.A(_14730_),
    .B1(_14805_),
    .B2(_15084_),
    .ZN(_15160_));
 NOR4_X1 _24871_ (.A1(_15157_),
    .A2(_15158_),
    .A3(_15159_),
    .A4(_15160_),
    .ZN(_15161_));
 NAND2_X1 _24872_ (.A1(_14755_),
    .A2(_14705_),
    .ZN(_15162_));
 OAI21_X1 _24873_ (.A(_14706_),
    .B1(_14988_),
    .B2(_14768_),
    .ZN(_15163_));
 AND4_X1 _24874_ (.A1(_14993_),
    .A2(_15161_),
    .A3(_15162_),
    .A4(_15163_),
    .ZN(_15164_));
 AOI21_X1 _24875_ (.A(_14946_),
    .B1(_14738_),
    .B2(_14880_),
    .ZN(_15165_));
 AND2_X1 _24876_ (.A1(_14752_),
    .A2(_14690_),
    .ZN(_15166_));
 INV_X1 _24877_ (.A(_15166_),
    .ZN(_15167_));
 NAND2_X1 _24878_ (.A1(_14761_),
    .A2(_14691_),
    .ZN(_15168_));
 OAI211_X1 _24879_ (.A(_14691_),
    .B(_14773_),
    .C1(_04132_),
    .C2(_09452_),
    .ZN(_15169_));
 NAND4_X1 _24880_ (.A1(_15167_),
    .A2(_14951_),
    .A3(_15168_),
    .A4(_15169_),
    .ZN(_15170_));
 NOR4_X1 _24881_ (.A1(_15165_),
    .A2(_15170_),
    .A3(_14841_),
    .A4(_14947_),
    .ZN(_15171_));
 NAND2_X1 _24882_ (.A1(_14883_),
    .A2(_14678_),
    .ZN(_15172_));
 NAND2_X1 _24883_ (.A1(_14883_),
    .A2(_14760_),
    .ZN(_15173_));
 OAI211_X1 _24884_ (.A(_15172_),
    .B(_15173_),
    .C1(_14667_),
    .C2(_14672_),
    .ZN(_15174_));
 OAI21_X1 _24885_ (.A(_14675_),
    .B1(_14901_),
    .B2(_14822_),
    .ZN(_15175_));
 OAI21_X1 _24886_ (.A(_15175_),
    .B1(_14811_),
    .B2(_14676_),
    .ZN(_15176_));
 AND2_X1 _24887_ (.A1(_14883_),
    .A2(_14714_),
    .ZN(_15177_));
 AND2_X1 _24888_ (.A1(_14883_),
    .A2(_14801_),
    .ZN(_15178_));
 NOR4_X1 _24889_ (.A1(_15174_),
    .A2(_15176_),
    .A3(_15177_),
    .A4(_15178_),
    .ZN(_15179_));
 NOR3_X1 _24890_ (.A1(_14712_),
    .A2(_17089_),
    .A3(_14699_),
    .ZN(_15180_));
 OAI21_X1 _24891_ (.A(_14717_),
    .B1(_14837_),
    .B2(_15180_),
    .ZN(_15181_));
 AND2_X1 _24892_ (.A1(_14821_),
    .A2(_14801_),
    .ZN(_15182_));
 AND2_X1 _24893_ (.A1(_14684_),
    .A2(_14748_),
    .ZN(_15183_));
 NOR4_X1 _24894_ (.A1(_15182_),
    .A2(_15112_),
    .A3(_15183_),
    .A4(_15111_),
    .ZN(_15184_));
 OAI21_X1 _24895_ (.A(_14821_),
    .B1(_14793_),
    .B2(_14924_),
    .ZN(_15185_));
 NAND2_X1 _24896_ (.A1(_14716_),
    .A2(_14681_),
    .ZN(_15186_));
 NAND2_X1 _24897_ (.A1(_14716_),
    .A2(_14671_),
    .ZN(_15187_));
 AND3_X1 _24898_ (.A1(_14829_),
    .A2(_15186_),
    .A3(_15187_),
    .ZN(_15188_));
 AND4_X1 _24899_ (.A1(_15181_),
    .A2(_15184_),
    .A3(_15185_),
    .A4(_15188_),
    .ZN(_15189_));
 NAND4_X1 _24900_ (.A1(_15164_),
    .A2(_15171_),
    .A3(_15179_),
    .A4(_15189_),
    .ZN(_15190_));
 AND2_X1 _24901_ (.A1(_14698_),
    .A2(_14761_),
    .ZN(_15191_));
 OR4_X1 _24902_ (.A1(_14910_),
    .A2(_15086_),
    .A3(_15191_),
    .A4(_15087_),
    .ZN(_15192_));
 AOI21_X1 _24903_ (.A(_14917_),
    .B1(_14940_),
    .B2(_14679_),
    .ZN(_15193_));
 NAND2_X1 _24904_ (.A1(_14781_),
    .A2(_14782_),
    .ZN(_15194_));
 OAI221_X1 _24905_ (.A(_15194_),
    .B1(_14913_),
    .B2(_14679_),
    .C1(_15028_),
    .C2(_04132_),
    .ZN(_15195_));
 NOR4_X1 _24906_ (.A1(_15192_),
    .A2(_15024_),
    .A3(_15193_),
    .A4(_15195_),
    .ZN(_15196_));
 AOI21_X1 _24907_ (.A(_14962_),
    .B1(_14790_),
    .B2(_15103_),
    .ZN(_15197_));
 AOI21_X1 _24908_ (.A(_14962_),
    .B1(_14899_),
    .B2(_14987_),
    .ZN(_15198_));
 AOI21_X1 _24909_ (.A(_15038_),
    .B1(_14710_),
    .B2(_14899_),
    .ZN(_15199_));
 NOR4_X1 _24910_ (.A1(_15197_),
    .A2(_15198_),
    .A3(_15199_),
    .A4(_14967_),
    .ZN(_15200_));
 AND2_X1 _24911_ (.A1(_14866_),
    .A2(_14869_),
    .ZN(_15201_));
 AND2_X1 _24912_ (.A1(_14826_),
    .A2(_14782_),
    .ZN(_15202_));
 NOR3_X1 _24913_ (.A1(_14972_),
    .A2(_15070_),
    .A3(_15202_),
    .ZN(_15203_));
 OAI21_X1 _24914_ (.A(_14956_),
    .B1(_14760_),
    .B2(_14782_),
    .ZN(_15204_));
 OAI21_X1 _24915_ (.A(_14956_),
    .B1(_14906_),
    .B2(_14984_),
    .ZN(_15205_));
 AND4_X1 _24916_ (.A1(_15201_),
    .A2(_15203_),
    .A3(_15204_),
    .A4(_15205_),
    .ZN(_15206_));
 INV_X1 _24917_ (.A(_15094_),
    .ZN(_15207_));
 OAI211_X1 _24918_ (.A(_15207_),
    .B(_15096_),
    .C1(_14810_),
    .C2(_14880_),
    .ZN(_15208_));
 AOI21_X1 _24919_ (.A(_14806_),
    .B1(_14916_),
    .B2(_14895_),
    .ZN(_15209_));
 NOR4_X1 _24920_ (.A1(_15208_),
    .A2(_15058_),
    .A3(_14922_),
    .A4(_15209_),
    .ZN(_15210_));
 NAND4_X1 _24921_ (.A1(_15196_),
    .A2(_15200_),
    .A3(_15206_),
    .A4(_15210_),
    .ZN(_15211_));
 NOR2_X1 _24922_ (.A1(_15190_),
    .A2(_15211_),
    .ZN(_15212_));
 XOR2_X1 _24923_ (.A(_15212_),
    .B(_01001_),
    .Z(_15213_));
 MUX2_X1 _24924_ (.A(_01211_),
    .B(_15213_),
    .S(_15147_),
    .Z(_01061_));
 INV_X1 _24925_ (.A(_15086_),
    .ZN(_15214_));
 OAI21_X1 _24926_ (.A(_15214_),
    .B1(_14913_),
    .B2(_15010_),
    .ZN(_15215_));
 AND2_X1 _24927_ (.A1(_14698_),
    .A2(_14763_),
    .ZN(_15216_));
 AND2_X1 _24928_ (.A1(_14698_),
    .A2(_14678_),
    .ZN(_15217_));
 AND2_X1 _24929_ (.A1(_14698_),
    .A2(_14924_),
    .ZN(_15218_));
 NOR4_X1 _24930_ (.A1(_15215_),
    .A2(_15216_),
    .A3(_15217_),
    .A4(_15218_),
    .ZN(_15219_));
 AOI21_X1 _24931_ (.A(_15032_),
    .B1(_14678_),
    .B2(_14703_),
    .ZN(_15220_));
 NAND4_X1 _24932_ (.A1(_14703_),
    .A2(_14773_),
    .A3(_14708_),
    .A4(_14739_),
    .ZN(_15221_));
 OAI21_X1 _24933_ (.A(_14703_),
    .B1(_14984_),
    .B2(_15115_),
    .ZN(_15222_));
 NAND4_X1 _24934_ (.A1(_15219_),
    .A2(_15220_),
    .A3(_15221_),
    .A4(_15222_),
    .ZN(_15223_));
 AND3_X1 _24935_ (.A1(_14789_),
    .A2(_14867_),
    .A3(_14673_),
    .ZN(_15224_));
 OAI211_X1 _24936_ (.A(_14831_),
    .B(_14701_),
    .C1(_17067_),
    .C2(_09041_),
    .ZN(_15225_));
 OAI21_X1 _24937_ (.A(_14831_),
    .B1(_14752_),
    .B2(_14747_),
    .ZN(_15226_));
 NAND2_X1 _24938_ (.A1(_15225_),
    .A2(_15226_),
    .ZN(_15227_));
 AOI21_X1 _24939_ (.A(_14962_),
    .B1(_14805_),
    .B2(_14792_),
    .ZN(_15228_));
 OR4_X1 _24940_ (.A1(_15224_),
    .A2(_15080_),
    .A3(_15227_),
    .A4(_15228_),
    .ZN(_15229_));
 AND2_X1 _24941_ (.A1(_14826_),
    .A2(_14744_),
    .ZN(_15230_));
 AOI211_X1 _24942_ (.A(_15230_),
    .B(_15067_),
    .C1(_14857_),
    .C2(_14865_),
    .ZN(_15231_));
 AND2_X1 _24943_ (.A1(_14800_),
    .A2(_14816_),
    .ZN(_15232_));
 AND2_X1 _24944_ (.A1(_14768_),
    .A2(_14816_),
    .ZN(_15233_));
 AND2_X1 _24945_ (.A1(_14815_),
    .A2(_14714_),
    .ZN(_15234_));
 AND2_X1 _24946_ (.A1(_14815_),
    .A2(_14687_),
    .ZN(_15235_));
 NOR4_X1 _24947_ (.A1(_15232_),
    .A2(_15233_),
    .A3(_15234_),
    .A4(_15235_),
    .ZN(_15236_));
 NAND2_X1 _24948_ (.A1(_14826_),
    .A2(_14777_),
    .ZN(_15237_));
 INV_X1 _24949_ (.A(_15202_),
    .ZN(_15238_));
 NAND2_X1 _24950_ (.A1(_14924_),
    .A2(_14826_),
    .ZN(_15239_));
 NAND3_X1 _24951_ (.A1(_14796_),
    .A2(_14749_),
    .A3(_14723_),
    .ZN(_15240_));
 AND4_X1 _24952_ (.A1(_15237_),
    .A2(_15238_),
    .A3(_15239_),
    .A4(_15240_),
    .ZN(_15241_));
 OAI21_X1 _24953_ (.A(_14956_),
    .B1(_14888_),
    .B2(_14819_),
    .ZN(_15242_));
 NAND4_X1 _24954_ (.A1(_15231_),
    .A2(_15236_),
    .A3(_15241_),
    .A4(_15242_),
    .ZN(_15243_));
 NOR3_X1 _24955_ (.A1(_14780_),
    .A2(_15097_),
    .A3(_14930_),
    .ZN(_15244_));
 OAI21_X1 _24956_ (.A(_14788_),
    .B1(_14801_),
    .B2(_14857_),
    .ZN(_15245_));
 OAI21_X1 _24957_ (.A(_14788_),
    .B1(_14755_),
    .B2(_14678_),
    .ZN(_15246_));
 OAI21_X1 _24958_ (.A(_14779_),
    .B1(_14892_),
    .B2(_15135_),
    .ZN(_15247_));
 NAND4_X1 _24959_ (.A1(_15244_),
    .A2(_15245_),
    .A3(_15246_),
    .A4(_15247_),
    .ZN(_15248_));
 NOR4_X1 _24960_ (.A1(_15223_),
    .A2(_15229_),
    .A3(_15243_),
    .A4(_15248_),
    .ZN(_15249_));
 NAND2_X1 _24961_ (.A1(_14756_),
    .A2(_15084_),
    .ZN(_15250_));
 AND2_X1 _24962_ (.A1(_15250_),
    .A2(_14942_),
    .ZN(_15251_));
 AND3_X1 _24963_ (.A1(_14808_),
    .A2(_14942_),
    .A3(_14739_),
    .ZN(_15252_));
 AOI21_X1 _24964_ (.A(_14730_),
    .B1(_15012_),
    .B2(_14899_),
    .ZN(_15253_));
 OR4_X1 _24965_ (.A1(_15158_),
    .A2(_15251_),
    .A3(_15252_),
    .A4(_15253_),
    .ZN(_15254_));
 NOR2_X1 _24966_ (.A1(_14766_),
    .A2(_14740_),
    .ZN(_15255_));
 AOI221_X4 _24967_ (.A(_14766_),
    .B1(_04121_),
    .B2(_09452_),
    .C1(_14880_),
    .C2(_14811_),
    .ZN(_15256_));
 NOR4_X1 _24968_ (.A1(_15254_),
    .A2(_14994_),
    .A3(_15255_),
    .A4(_15256_),
    .ZN(_15257_));
 AND2_X1 _24969_ (.A1(_14856_),
    .A2(_14690_),
    .ZN(_15258_));
 INV_X1 _24970_ (.A(_15258_),
    .ZN(_15259_));
 NAND4_X1 _24971_ (.A1(_15259_),
    .A2(_15167_),
    .A3(_14949_),
    .A4(_14951_),
    .ZN(_15260_));
 OAI211_X1 _24972_ (.A(_15003_),
    .B(_15005_),
    .C1(_14740_),
    .C2(_14946_),
    .ZN(_15261_));
 NAND2_X1 _24973_ (.A1(_14751_),
    .A2(_14714_),
    .ZN(_15262_));
 NAND4_X1 _24974_ (.A1(_14749_),
    .A2(_14783_),
    .A3(_14837_),
    .A4(_14764_),
    .ZN(_15263_));
 OAI211_X1 _24975_ (.A(_15262_),
    .B(_15263_),
    .C1(_15010_),
    .C2(_14946_),
    .ZN(_15264_));
 AND4_X1 _24976_ (.A1(_14858_),
    .A2(_14732_),
    .A3(_14764_),
    .A4(_14770_),
    .ZN(_15265_));
 NOR4_X1 _24977_ (.A1(_15260_),
    .A2(_15261_),
    .A3(_15264_),
    .A4(_15265_),
    .ZN(_15266_));
 OAI21_X1 _24978_ (.A(_14675_),
    .B1(_14782_),
    .B2(_14719_),
    .ZN(_15267_));
 AND3_X1 _24979_ (.A1(_15267_),
    .A2(_14802_),
    .A3(_14804_),
    .ZN(_15268_));
 NAND3_X1 _24980_ (.A1(_14924_),
    .A2(_14665_),
    .A3(_14803_),
    .ZN(_15269_));
 OAI21_X1 _24981_ (.A(_15269_),
    .B1(_14667_),
    .B2(_14805_),
    .ZN(_15270_));
 AND2_X1 _24982_ (.A1(_14883_),
    .A2(_14789_),
    .ZN(_15271_));
 AND4_X1 _24983_ (.A1(_14707_),
    .A2(_14662_),
    .A3(_14665_),
    .A4(_14701_),
    .ZN(_15272_));
 NOR4_X1 _24984_ (.A1(_15270_),
    .A2(_15271_),
    .A3(_15177_),
    .A4(_15272_),
    .ZN(_15273_));
 NAND2_X1 _24985_ (.A1(_14684_),
    .A2(_14702_),
    .ZN(_15274_));
 OAI21_X1 _24986_ (.A(_15274_),
    .B1(_14757_),
    .B2(_15013_),
    .ZN(_15275_));
 AND2_X1 _24987_ (.A1(_14684_),
    .A2(_14924_),
    .ZN(_15276_));
 NOR3_X1 _24988_ (.A1(_15275_),
    .A2(_15276_),
    .A3(_14897_),
    .ZN(_15277_));
 NAND2_X1 _24989_ (.A1(_14717_),
    .A2(_14777_),
    .ZN(_15278_));
 OAI21_X1 _24990_ (.A(_14716_),
    .B1(_14857_),
    .B2(_14884_),
    .ZN(_15279_));
 AND4_X1 _24991_ (.A1(_15278_),
    .A2(_14855_),
    .A3(_15279_),
    .A4(_15187_),
    .ZN(_15280_));
 AND4_X1 _24992_ (.A1(_15268_),
    .A2(_15273_),
    .A3(_15277_),
    .A4(_15280_),
    .ZN(_15281_));
 NAND4_X1 _24993_ (.A1(_15249_),
    .A2(_15257_),
    .A3(_15266_),
    .A4(_15281_),
    .ZN(_15282_));
 NOR2_X1 _24994_ (.A1(_15282_),
    .A2(_14797_),
    .ZN(_15283_));
 INV_X1 _24995_ (.A(_01002_),
    .ZN(_15284_));
 XNOR2_X1 _24996_ (.A(_15283_),
    .B(_15284_),
    .ZN(_15285_));
 MUX2_X1 _24997_ (.A(_01212_),
    .B(_15285_),
    .S(_15147_),
    .Z(_01062_));
 OR2_X1 _24998_ (.A1(_14827_),
    .A2(_15070_),
    .ZN(_15286_));
 AND3_X1 _24999_ (.A1(_14796_),
    .A2(_14749_),
    .A3(_14867_),
    .ZN(_15287_));
 OR4_X1 _25000_ (.A1(_15230_),
    .A2(_15286_),
    .A3(_14971_),
    .A4(_15287_),
    .ZN(_15288_));
 OAI21_X1 _25001_ (.A(_14832_),
    .B1(_14793_),
    .B2(_14901_),
    .ZN(_15289_));
 NAND2_X1 _25002_ (.A1(_14832_),
    .A2(_14753_),
    .ZN(_15290_));
 NAND4_X1 _25003_ (.A1(_14851_),
    .A2(_14867_),
    .A3(_14783_),
    .A4(_14673_),
    .ZN(_15291_));
 NAND4_X1 _25004_ (.A1(_15289_),
    .A2(_15290_),
    .A3(_15040_),
    .A4(_15291_),
    .ZN(_15292_));
 NAND2_X1 _25005_ (.A1(_14988_),
    .A2(_14725_),
    .ZN(_15293_));
 OAI211_X1 _25006_ (.A(_14850_),
    .B(_14867_),
    .C1(_14796_),
    .C2(_14763_),
    .ZN(_15294_));
 OAI211_X1 _25007_ (.A(_15293_),
    .B(_15294_),
    .C1(_15010_),
    .C2(_14962_),
    .ZN(_15295_));
 OAI21_X1 _25008_ (.A(_14956_),
    .B1(_14822_),
    .B2(_14678_),
    .ZN(_15296_));
 OAI211_X1 _25009_ (.A(_14956_),
    .B(_17092_),
    .C1(_09452_),
    .C2(_14668_),
    .ZN(_15297_));
 INV_X1 _25010_ (.A(_14956_),
    .ZN(_15298_));
 OAI211_X1 _25011_ (.A(_15296_),
    .B(_15297_),
    .C1(_14742_),
    .C2(_15298_),
    .ZN(_15299_));
 NOR4_X1 _25012_ (.A1(_15288_),
    .A2(_15292_),
    .A3(_15295_),
    .A4(_15299_),
    .ZN(_15300_));
 OAI21_X1 _25013_ (.A(_14942_),
    .B1(_14819_),
    .B2(_14773_),
    .ZN(_15301_));
 AND2_X1 _25014_ (.A1(_14747_),
    .A2(_14690_),
    .ZN(_15302_));
 AND2_X1 _25015_ (.A1(_14690_),
    .A2(_14720_),
    .ZN(_15303_));
 NOR4_X1 _25016_ (.A1(_15166_),
    .A2(_15258_),
    .A3(_15302_),
    .A4(_15303_),
    .ZN(_15304_));
 OAI21_X1 _25017_ (.A(_14750_),
    .B1(_14984_),
    .B2(_14748_),
    .ZN(_15305_));
 OAI21_X1 _25018_ (.A(_14750_),
    .B1(_14777_),
    .B2(_14671_),
    .ZN(_15306_));
 AND4_X1 _25019_ (.A1(_15262_),
    .A2(_15304_),
    .A3(_15305_),
    .A4(_15306_),
    .ZN(_15307_));
 NAND3_X1 _25020_ (.A1(_14705_),
    .A2(_14718_),
    .A3(_14735_),
    .ZN(_15308_));
 OAI211_X1 _25021_ (.A(_15162_),
    .B(_15308_),
    .C1(_14672_),
    .C2(_14766_),
    .ZN(_15309_));
 AND3_X1 _25022_ (.A1(_14705_),
    .A2(_14732_),
    .A3(_14701_),
    .ZN(_15310_));
 NOR2_X1 _25023_ (.A1(_14766_),
    .A2(_14987_),
    .ZN(_15311_));
 NOR4_X1 _25024_ (.A1(_15309_),
    .A2(_14994_),
    .A3(_15310_),
    .A4(_15311_),
    .ZN(_15312_));
 AOI211_X1 _25025_ (.A(_14943_),
    .B(_15159_),
    .C1(_14942_),
    .C2(_14753_),
    .ZN(_15313_));
 AND4_X1 _25026_ (.A1(_15301_),
    .A2(_15307_),
    .A3(_15312_),
    .A4(_15313_),
    .ZN(_15314_));
 AND2_X1 _25027_ (.A1(_14683_),
    .A2(_14763_),
    .ZN(_15315_));
 AOI221_X4 _25028_ (.A(_14981_),
    .B1(_14681_),
    .B2(_14684_),
    .C1(_04121_),
    .C2(_15315_),
    .ZN(_15316_));
 NAND2_X1 _25029_ (.A1(_14821_),
    .A2(_14748_),
    .ZN(_15317_));
 NAND3_X1 _25030_ (.A1(_15316_),
    .A2(_14846_),
    .A3(_15317_),
    .ZN(_15318_));
 NOR2_X1 _25031_ (.A1(_15139_),
    .A2(_14885_),
    .ZN(_15319_));
 OAI211_X1 _25032_ (.A(_15319_),
    .B(_15141_),
    .C1(_14861_),
    .C2(_14667_),
    .ZN(_15320_));
 OAI21_X1 _25033_ (.A(_14675_),
    .B1(_14984_),
    .B2(_15115_),
    .ZN(_15321_));
 OAI21_X1 _25034_ (.A(_15321_),
    .B1(_14742_),
    .B2(_14676_),
    .ZN(_15322_));
 AND2_X1 _25035_ (.A1(_14716_),
    .A2(_14872_),
    .ZN(_15323_));
 AND2_X1 _25036_ (.A1(_14716_),
    .A2(_14891_),
    .ZN(_15324_));
 AND3_X1 _25037_ (.A1(_14888_),
    .A2(_14858_),
    .A3(_14662_),
    .ZN(_15325_));
 OR4_X1 _25038_ (.A1(_15323_),
    .A2(_14903_),
    .A3(_15324_),
    .A4(_15325_),
    .ZN(_15326_));
 NOR4_X1 _25039_ (.A1(_15318_),
    .A2(_15320_),
    .A3(_15322_),
    .A4(_15326_),
    .ZN(_15327_));
 OAI21_X1 _25040_ (.A(_14781_),
    .B1(_14984_),
    .B2(_15115_),
    .ZN(_15328_));
 OAI211_X1 _25041_ (.A(_14694_),
    .B(_14665_),
    .C1(_14789_),
    .C2(_14796_),
    .ZN(_15329_));
 NAND4_X1 _25042_ (.A1(_14850_),
    .A2(_14783_),
    .A3(_14773_),
    .A4(_14694_),
    .ZN(_15330_));
 AND3_X1 _25043_ (.A1(_15328_),
    .A2(_15329_),
    .A3(_15330_),
    .ZN(_15331_));
 INV_X1 _25044_ (.A(_15060_),
    .ZN(_15332_));
 AND2_X1 _25045_ (.A1(_14787_),
    .A2(_14857_),
    .ZN(_15333_));
 AND2_X1 _25046_ (.A1(_14681_),
    .A2(_14787_),
    .ZN(_15334_));
 AND2_X1 _25047_ (.A1(_14787_),
    .A2(_14678_),
    .ZN(_15335_));
 NOR4_X1 _25048_ (.A1(_15332_),
    .A2(_15333_),
    .A3(_15334_),
    .A4(_15335_),
    .ZN(_15336_));
 AOI21_X1 _25049_ (.A(_14917_),
    .B1(_15101_),
    .B2(_15084_),
    .ZN(_15337_));
 AND2_X1 _25050_ (.A1(_14892_),
    .A2(_14703_),
    .ZN(_15338_));
 NOR4_X1 _25051_ (.A1(_15337_),
    .A2(_15338_),
    .A3(_15090_),
    .A4(_14920_),
    .ZN(_15339_));
 OAI21_X1 _25052_ (.A(_14779_),
    .B1(_14854_),
    .B2(_14768_),
    .ZN(_15340_));
 NAND3_X1 _25053_ (.A1(_14779_),
    .A2(_14718_),
    .A3(_14735_),
    .ZN(_15341_));
 AND4_X1 _25054_ (.A1(_14934_),
    .A2(_15098_),
    .A3(_15340_),
    .A4(_15341_),
    .ZN(_15342_));
 AND4_X1 _25055_ (.A1(_15331_),
    .A2(_15336_),
    .A3(_15339_),
    .A4(_15342_),
    .ZN(_15343_));
 NAND4_X1 _25056_ (.A1(_15300_),
    .A2(_15314_),
    .A3(_15327_),
    .A4(_15343_),
    .ZN(_15344_));
 NOR2_X1 _25057_ (.A1(_15344_),
    .A2(_14797_),
    .ZN(_15345_));
 INV_X1 _25058_ (.A(_01003_),
    .ZN(_15346_));
 XNOR2_X1 _25059_ (.A(_15345_),
    .B(_15346_),
    .ZN(_15347_));
 MUX2_X1 _25060_ (.A(_01214_),
    .B(_15347_),
    .S(_15147_),
    .Z(_01063_));
 AND2_X1 _25061_ (.A1(_14942_),
    .A2(_14768_),
    .ZN(_15348_));
 AOI211_X1 _25062_ (.A(_14880_),
    .B(_14730_),
    .C1(_14734_),
    .C2(_09041_),
    .ZN(_15349_));
 OR4_X1 _25063_ (.A1(_15348_),
    .A2(_15349_),
    .A3(_14944_),
    .A4(_15159_),
    .ZN(_15350_));
 OAI21_X1 _25064_ (.A(_14706_),
    .B1(_14755_),
    .B2(_14888_),
    .ZN(_15351_));
 NAND3_X1 _25065_ (.A1(_15351_),
    .A2(_15126_),
    .A3(_15124_),
    .ZN(_15352_));
 AOI21_X1 _25066_ (.A(_14730_),
    .B1(_15031_),
    .B2(_14679_),
    .ZN(_15353_));
 NOR4_X1 _25067_ (.A1(_15350_),
    .A2(_15352_),
    .A3(_15251_),
    .A4(_15353_),
    .ZN(_15354_));
 NAND2_X1 _25068_ (.A1(_14683_),
    .A2(_14761_),
    .ZN(_15355_));
 OAI21_X1 _25069_ (.A(_15355_),
    .B1(_14757_),
    .B2(_15156_),
    .ZN(_15356_));
 OR4_X1 _25070_ (.A1(_14980_),
    .A2(_15356_),
    .A3(_15315_),
    .A4(_14981_),
    .ZN(_15357_));
 AND2_X1 _25071_ (.A1(_14717_),
    .A2(_15180_),
    .ZN(_15358_));
 NAND3_X1 _25072_ (.A1(_14888_),
    .A2(_14858_),
    .A3(_14803_),
    .ZN(_15359_));
 OAI211_X1 _25073_ (.A(_15186_),
    .B(_15359_),
    .C1(_14904_),
    .C2(_14878_),
    .ZN(_15360_));
 NOR4_X1 _25074_ (.A1(_15357_),
    .A2(_14903_),
    .A3(_15358_),
    .A4(_15360_),
    .ZN(_15361_));
 NAND4_X1 _25075_ (.A1(_14842_),
    .A2(_14844_),
    .A3(_15006_),
    .A4(_15129_),
    .ZN(_15362_));
 AND4_X1 _25076_ (.A1(_09041_),
    .A2(_14851_),
    .A3(_14858_),
    .A4(_14764_),
    .ZN(_15363_));
 NAND2_X1 _25077_ (.A1(_14951_),
    .A2(_15132_),
    .ZN(_15364_));
 AOI21_X1 _25078_ (.A(_15001_),
    .B1(_14916_),
    .B2(_14878_),
    .ZN(_15365_));
 NOR4_X1 _25079_ (.A1(_15362_),
    .A2(_15363_),
    .A3(_15364_),
    .A4(_15365_),
    .ZN(_15366_));
 OAI211_X1 _25080_ (.A(_15173_),
    .B(_15269_),
    .C1(_14667_),
    .C2(_14878_),
    .ZN(_15367_));
 AOI21_X1 _25081_ (.A(_14676_),
    .B1(_15101_),
    .B2(_15084_),
    .ZN(_15368_));
 AOI21_X1 _25082_ (.A(_14676_),
    .B1(_15013_),
    .B2(_14899_),
    .ZN(_15369_));
 NAND3_X1 _25083_ (.A1(_14883_),
    .A2(_14843_),
    .A3(_14739_),
    .ZN(_15370_));
 NAND2_X1 _25084_ (.A1(_15370_),
    .A2(_14849_),
    .ZN(_15371_));
 NOR4_X1 _25085_ (.A1(_15367_),
    .A2(_15368_),
    .A3(_15369_),
    .A4(_15371_),
    .ZN(_15372_));
 AND4_X1 _25086_ (.A1(_15354_),
    .A2(_15361_),
    .A3(_15366_),
    .A4(_15372_),
    .ZN(_15373_));
 AND2_X1 _25087_ (.A1(_14884_),
    .A2(_14831_),
    .ZN(_15374_));
 INV_X1 _25088_ (.A(_15374_),
    .ZN(_15375_));
 NOR2_X1 _25089_ (.A1(_14752_),
    .A2(_14747_),
    .ZN(_15376_));
 NOR2_X1 _25090_ (.A1(_14962_),
    .A2(_15376_),
    .ZN(_15377_));
 AOI21_X1 _25091_ (.A(_15377_),
    .B1(_14725_),
    .B2(_14906_),
    .ZN(_15378_));
 OAI21_X1 _25092_ (.A(_14725_),
    .B1(_14671_),
    .B2(_14720_),
    .ZN(_15379_));
 OAI21_X1 _25093_ (.A(_14831_),
    .B1(_14793_),
    .B2(_14760_),
    .ZN(_15380_));
 AND4_X1 _25094_ (.A1(_15375_),
    .A2(_15378_),
    .A3(_15379_),
    .A4(_15380_),
    .ZN(_15381_));
 AND2_X1 _25095_ (.A1(_14727_),
    .A2(_14778_),
    .ZN(_15382_));
 AND2_X1 _25096_ (.A1(_14778_),
    .A2(_15135_),
    .ZN(_15383_));
 OR4_X1 _25097_ (.A1(_14930_),
    .A2(_15094_),
    .A3(_15382_),
    .A4(_15383_),
    .ZN(_15384_));
 AOI21_X1 _25098_ (.A(_14806_),
    .B1(_15031_),
    .B2(_14679_),
    .ZN(_15385_));
 NAND2_X1 _25099_ (.A1(_14760_),
    .A2(_14788_),
    .ZN(_15386_));
 NAND2_X1 _25100_ (.A1(_15386_),
    .A2(_15053_),
    .ZN(_15387_));
 NAND2_X1 _25101_ (.A1(_14928_),
    .A2(_14864_),
    .ZN(_15388_));
 NOR4_X1 _25102_ (.A1(_15384_),
    .A2(_15385_),
    .A3(_15387_),
    .A4(_15388_),
    .ZN(_15389_));
 NOR2_X1 _25103_ (.A1(_15232_),
    .A2(_15234_),
    .ZN(_15390_));
 AND2_X1 _25104_ (.A1(_14815_),
    .A2(_14678_),
    .ZN(_15391_));
 AND2_X1 _25105_ (.A1(_14815_),
    .A2(_14888_),
    .ZN(_15392_));
 AOI211_X1 _25106_ (.A(_15391_),
    .B(_15392_),
    .C1(_14681_),
    .C2(_14816_),
    .ZN(_15393_));
 OAI221_X1 _25107_ (.A(_14865_),
    .B1(_14734_),
    .B2(_09452_),
    .C1(_14837_),
    .C2(_14851_),
    .ZN(_15394_));
 AND4_X1 _25108_ (.A1(_15390_),
    .A2(_15393_),
    .A3(_15240_),
    .A4(_15394_),
    .ZN(_15395_));
 INV_X1 _25109_ (.A(_15218_),
    .ZN(_15396_));
 OAI211_X1 _25110_ (.A(_14694_),
    .B(_14665_),
    .C1(_14753_),
    .C2(_14687_),
    .ZN(_15397_));
 NAND4_X1 _25111_ (.A1(_15214_),
    .A2(_15396_),
    .A3(_15194_),
    .A4(_15397_),
    .ZN(_15398_));
 AND2_X1 _25112_ (.A1(_14703_),
    .A2(_14796_),
    .ZN(_15399_));
 AND2_X1 _25113_ (.A1(_15030_),
    .A2(_14708_),
    .ZN(_15400_));
 OAI211_X1 _25114_ (.A(_14695_),
    .B(_14837_),
    .C1(_04121_),
    .C2(_09041_),
    .ZN(_15401_));
 OAI21_X1 _25115_ (.A(_15401_),
    .B1(_15010_),
    .B2(_14917_),
    .ZN(_15402_));
 NOR4_X1 _25116_ (.A1(_15398_),
    .A2(_15399_),
    .A3(_15400_),
    .A4(_15402_),
    .ZN(_15403_));
 AND4_X1 _25117_ (.A1(_15381_),
    .A2(_15389_),
    .A3(_15395_),
    .A4(_15403_),
    .ZN(_15404_));
 AND2_X1 _25118_ (.A1(_15373_),
    .A2(_15404_),
    .ZN(_15405_));
 INV_X1 _25119_ (.A(_01004_),
    .ZN(_15406_));
 XNOR2_X1 _25120_ (.A(_15405_),
    .B(_15406_),
    .ZN(_15407_));
 MUX2_X1 _25121_ (.A(_01215_),
    .B(_15407_),
    .S(_15147_),
    .Z(_01064_));
 NOR2_X1 _25122_ (.A1(_10970_),
    .A2(_17070_),
    .ZN(_15408_));
 CLKBUF_X2 _25123_ (.A(_15408_),
    .Z(_15409_));
 NOR2_X1 _25124_ (.A1(_10976_),
    .A2(_17073_),
    .ZN(_15410_));
 AND2_X1 _25125_ (.A1(_15409_),
    .A2(_15410_),
    .ZN(_15411_));
 CLKBUF_X2 _25126_ (.A(_15411_),
    .Z(_15412_));
 BUF_X2 _25127_ (.A(_15412_),
    .Z(_15413_));
 AND2_X1 _25128_ (.A1(_10931_),
    .A2(_17098_),
    .ZN(_15414_));
 CLKBUF_X2 _25129_ (.A(_15414_),
    .Z(_15415_));
 NOR2_X1 _25130_ (.A1(_17068_),
    .A2(_17069_),
    .ZN(_15416_));
 CLKBUF_X2 _25131_ (.A(_15416_),
    .Z(_15417_));
 AND2_X1 _25132_ (.A1(_15415_),
    .A2(_15417_),
    .ZN(_15418_));
 CLKBUF_X2 _25133_ (.A(_15418_),
    .Z(_15419_));
 AND2_X1 _25134_ (.A1(_15413_),
    .A2(_15419_),
    .ZN(_15420_));
 INV_X1 _25135_ (.A(_15420_),
    .ZN(_15421_));
 INV_X1 _25136_ (.A(_17097_),
    .ZN(_15422_));
 NOR2_X1 _25137_ (.A1(_15422_),
    .A2(_17098_),
    .ZN(_15423_));
 CLKBUF_X2 _25138_ (.A(_15423_),
    .Z(_15424_));
 AND2_X1 _25139_ (.A1(_15424_),
    .A2(_15417_),
    .ZN(_15425_));
 AND2_X1 _25140_ (.A1(_15412_),
    .A2(_15425_),
    .ZN(_15426_));
 INV_X1 _25141_ (.A(_15426_),
    .ZN(_15427_));
 AND2_X1 _25142_ (.A1(_17070_),
    .A2(_17071_),
    .ZN(_15428_));
 CLKBUF_X2 _25143_ (.A(_15428_),
    .Z(_15429_));
 AND2_X2 _25144_ (.A1(_15410_),
    .A2(_15429_),
    .ZN(_15430_));
 CLKBUF_X2 _25145_ (.A(_15430_),
    .Z(_15431_));
 NOR2_X1 _25146_ (.A1(_10931_),
    .A2(_17098_),
    .ZN(_15432_));
 AND2_X1 _25147_ (.A1(_15432_),
    .A2(_15417_),
    .ZN(_15433_));
 BUF_X2 _25148_ (.A(_15433_),
    .Z(_15434_));
 NAND2_X1 _25149_ (.A1(_15431_),
    .A2(_15434_),
    .ZN(_15435_));
 CLKBUF_X2 _25150_ (.A(_15422_),
    .Z(_15436_));
 BUF_X2 _25151_ (.A(_15436_),
    .Z(_15437_));
 AND2_X1 _25152_ (.A1(_17068_),
    .A2(_17069_),
    .ZN(_15438_));
 AND2_X1 _25153_ (.A1(_15438_),
    .A2(_17098_),
    .ZN(_15439_));
 CLKBUF_X2 _25154_ (.A(_15439_),
    .Z(_15440_));
 NAND3_X1 _25155_ (.A1(_15413_),
    .A2(_15437_),
    .A3(_15440_),
    .ZN(_15441_));
 NAND4_X1 _25156_ (.A1(_15421_),
    .A2(_15427_),
    .A3(_15435_),
    .A4(_15441_),
    .ZN(_15442_));
 NOR2_X2 _25157_ (.A1(_17072_),
    .A2(_17073_),
    .ZN(_15443_));
 AND2_X1 _25158_ (.A1(_15409_),
    .A2(_15443_),
    .ZN(_15444_));
 CLKBUF_X2 _25159_ (.A(_15444_),
    .Z(_15445_));
 INV_X1 _25160_ (.A(_15417_),
    .ZN(_15446_));
 NOR2_X1 _25161_ (.A1(_15446_),
    .A2(_15415_),
    .ZN(_15447_));
 AND2_X1 _25162_ (.A1(_15445_),
    .A2(_15447_),
    .ZN(_15448_));
 NOR2_X2 _25163_ (.A1(_10964_),
    .A2(_17071_),
    .ZN(_15449_));
 AND2_X1 _25164_ (.A1(_17072_),
    .A2(_17073_),
    .ZN(_15450_));
 CLKBUF_X2 _25165_ (.A(_15450_),
    .Z(_15451_));
 AND2_X1 _25166_ (.A1(_15449_),
    .A2(_15451_),
    .ZN(_15452_));
 CLKBUF_X2 _25167_ (.A(_15452_),
    .Z(_15453_));
 INV_X1 _25168_ (.A(_17068_),
    .ZN(_15454_));
 NAND2_X1 _25169_ (.A1(_15454_),
    .A2(_17098_),
    .ZN(_15455_));
 NOR2_X2 _25170_ (.A1(_15455_),
    .A2(_17069_),
    .ZN(_15456_));
 AND2_X1 _25171_ (.A1(_15453_),
    .A2(_15456_),
    .ZN(_15457_));
 AND2_X1 _25172_ (.A1(_15457_),
    .A2(_15437_),
    .ZN(_15458_));
 BUF_X2 _25173_ (.A(_15432_),
    .Z(_15459_));
 INV_X1 _25174_ (.A(_15459_),
    .ZN(_15460_));
 INV_X1 _25175_ (.A(_17069_),
    .ZN(_15461_));
 NOR2_X1 _25176_ (.A1(_15461_),
    .A2(_17068_),
    .ZN(_15462_));
 CLKBUF_X2 _25177_ (.A(_15462_),
    .Z(_15463_));
 BUF_X2 _25178_ (.A(_15463_),
    .Z(_15464_));
 NAND2_X1 _25179_ (.A1(_15460_),
    .A2(_15464_),
    .ZN(_15465_));
 INV_X1 _25180_ (.A(_15409_),
    .ZN(_15466_));
 INV_X1 _25181_ (.A(_15443_),
    .ZN(_15467_));
 NOR3_X1 _25182_ (.A1(_15465_),
    .A2(_15466_),
    .A3(_15467_),
    .ZN(_15468_));
 NOR2_X2 _25183_ (.A1(_17070_),
    .A2(_17071_),
    .ZN(_15469_));
 AND2_X1 _25184_ (.A1(_15451_),
    .A2(_15469_),
    .ZN(_15470_));
 CLKBUF_X2 _25185_ (.A(_15470_),
    .Z(_15471_));
 CLKBUF_X2 _25186_ (.A(_15438_),
    .Z(_15472_));
 CLKBUF_X2 _25187_ (.A(_15472_),
    .Z(_15473_));
 NOR2_X1 _25188_ (.A1(_10944_),
    .A2(_10931_),
    .ZN(_15474_));
 CLKBUF_X2 _25189_ (.A(_15474_),
    .Z(_15475_));
 AND3_X1 _25190_ (.A1(_15471_),
    .A2(_15473_),
    .A3(_15475_),
    .ZN(_15476_));
 OR4_X1 _25191_ (.A1(_15448_),
    .A2(_15458_),
    .A3(_15468_),
    .A4(_15476_),
    .ZN(_15477_));
 NOR2_X2 _25192_ (.A1(_15454_),
    .A2(_17069_),
    .ZN(_15478_));
 AND2_X2 _25193_ (.A1(_15478_),
    .A2(_15432_),
    .ZN(_15479_));
 AND2_X1 _25194_ (.A1(_15428_),
    .A2(_15450_),
    .ZN(_15480_));
 AND2_X1 _25195_ (.A1(_15479_),
    .A2(_15480_),
    .ZN(_15481_));
 INV_X1 _25196_ (.A(_15481_),
    .ZN(_15482_));
 AND2_X1 _25197_ (.A1(_15408_),
    .A2(_15451_),
    .ZN(_15483_));
 CLKBUF_X2 _25198_ (.A(_15483_),
    .Z(_15484_));
 BUF_X2 _25199_ (.A(_15484_),
    .Z(_15485_));
 BUF_X2 _25200_ (.A(_15475_),
    .Z(_15486_));
 OAI211_X1 _25201_ (.A(_15485_),
    .B(_15464_),
    .C1(_15486_),
    .C2(_15415_),
    .ZN(_15487_));
 NAND4_X1 _25202_ (.A1(_15409_),
    .A2(_15464_),
    .A3(_15459_),
    .A4(_15451_),
    .ZN(_15488_));
 NAND2_X1 _25203_ (.A1(_15425_),
    .A2(_15480_),
    .ZN(_15489_));
 NAND4_X1 _25204_ (.A1(_15482_),
    .A2(_15487_),
    .A3(_15488_),
    .A4(_15489_),
    .ZN(_15490_));
 AND2_X1 _25205_ (.A1(_15424_),
    .A2(_15478_),
    .ZN(_15491_));
 AND2_X1 _25206_ (.A1(_15491_),
    .A2(_15453_),
    .ZN(_15492_));
 AND2_X2 _25207_ (.A1(_15474_),
    .A2(_15417_),
    .ZN(_15493_));
 AND2_X1 _25208_ (.A1(_15493_),
    .A2(_15470_),
    .ZN(_15494_));
 OR2_X1 _25209_ (.A1(_15492_),
    .A2(_15494_),
    .ZN(_15495_));
 NOR4_X1 _25210_ (.A1(_15442_),
    .A2(_15477_),
    .A3(_15490_),
    .A4(_15495_),
    .ZN(_15496_));
 AND2_X1 _25211_ (.A1(_15462_),
    .A2(_15432_),
    .ZN(_15497_));
 AND2_X2 _25212_ (.A1(_15429_),
    .A2(_15443_),
    .ZN(_15498_));
 CLKBUF_X2 _25213_ (.A(_15498_),
    .Z(_15499_));
 AND2_X1 _25214_ (.A1(_15497_),
    .A2(_15499_),
    .ZN(_15500_));
 NOR2_X1 _25215_ (.A1(_15446_),
    .A2(_15432_),
    .ZN(_15501_));
 AND2_X1 _25216_ (.A1(_15501_),
    .A2(_15499_),
    .ZN(_15502_));
 NOR2_X1 _25217_ (.A1(_15500_),
    .A2(_15502_),
    .ZN(_15503_));
 INV_X1 _25218_ (.A(_15438_),
    .ZN(_15504_));
 NOR2_X1 _25219_ (.A1(_15504_),
    .A2(_15459_),
    .ZN(_15505_));
 NOR2_X1 _25220_ (.A1(_10984_),
    .A2(_17072_),
    .ZN(_15506_));
 AND2_X1 _25221_ (.A1(_15506_),
    .A2(_15469_),
    .ZN(_15507_));
 AND2_X1 _25222_ (.A1(_15505_),
    .A2(_15507_),
    .ZN(_15508_));
 AND2_X1 _25223_ (.A1(_15506_),
    .A2(_15409_),
    .ZN(_15509_));
 AND2_X1 _25224_ (.A1(_15509_),
    .A2(_15479_),
    .ZN(_15510_));
 AND2_X1 _25225_ (.A1(_15506_),
    .A2(_15429_),
    .ZN(_15511_));
 BUF_X2 _25226_ (.A(_15511_),
    .Z(_15512_));
 BUF_X2 _25227_ (.A(_15512_),
    .Z(_15513_));
 NOR2_X1 _25228_ (.A1(_15446_),
    .A2(_15424_),
    .ZN(_15514_));
 AND2_X1 _25229_ (.A1(_15438_),
    .A2(_15432_),
    .ZN(_15515_));
 CLKBUF_X2 _25230_ (.A(_15515_),
    .Z(_15516_));
 NOR2_X1 _25231_ (.A1(_15514_),
    .A2(_15516_),
    .ZN(_15517_));
 INV_X1 _25232_ (.A(_15517_),
    .ZN(_15518_));
 AOI211_X1 _25233_ (.A(_15508_),
    .B(_15510_),
    .C1(_15513_),
    .C2(_15518_),
    .ZN(_15519_));
 AND2_X2 _25234_ (.A1(_15438_),
    .A2(_15415_),
    .ZN(_15520_));
 AND2_X1 _25235_ (.A1(_15520_),
    .A2(_15498_),
    .ZN(_15521_));
 AND2_X1 _25236_ (.A1(_15410_),
    .A2(_15469_),
    .ZN(_15522_));
 BUF_X2 _25237_ (.A(_15522_),
    .Z(_15523_));
 AND2_X2 _25238_ (.A1(_15478_),
    .A2(_17098_),
    .ZN(_15524_));
 AOI221_X4 _25239_ (.A(_15521_),
    .B1(_15479_),
    .B2(_15523_),
    .C1(_15524_),
    .C2(_15413_),
    .ZN(_15525_));
 AND2_X1 _25240_ (.A1(_15474_),
    .A2(_15478_),
    .ZN(_15526_));
 BUF_X2 _25241_ (.A(_15526_),
    .Z(_15527_));
 AOI22_X1 _25242_ (.A1(_15527_),
    .A2(_15499_),
    .B1(_15445_),
    .B2(_15516_),
    .ZN(_15528_));
 AND4_X1 _25243_ (.A1(_15503_),
    .A2(_15519_),
    .A3(_15525_),
    .A4(_15528_),
    .ZN(_15529_));
 AND2_X1 _25244_ (.A1(_15443_),
    .A2(_15469_),
    .ZN(_15530_));
 CLKBUF_X2 _25245_ (.A(_15530_),
    .Z(_15531_));
 CLKBUF_X2 _25246_ (.A(_15531_),
    .Z(_15532_));
 BUF_X2 _25247_ (.A(_15464_),
    .Z(_15533_));
 CLKBUF_X2 _25248_ (.A(_15478_),
    .Z(_15534_));
 CLKBUF_X2 _25249_ (.A(_15534_),
    .Z(_15535_));
 OAI211_X1 _25250_ (.A(_15532_),
    .B(_15424_),
    .C1(_15533_),
    .C2(_15535_),
    .ZN(_15536_));
 INV_X1 _25251_ (.A(_15456_),
    .ZN(_15537_));
 NAND3_X1 _25252_ (.A1(_10970_),
    .A2(_10976_),
    .A3(_10984_),
    .ZN(_15538_));
 INV_X1 _25253_ (.A(_15524_),
    .ZN(_15539_));
 INV_X1 _25254_ (.A(_15531_),
    .ZN(_15540_));
 OAI221_X1 _25255_ (.A(_15536_),
    .B1(_15537_),
    .B2(_15538_),
    .C1(_15539_),
    .C2(_15540_),
    .ZN(_15541_));
 AND2_X1 _25256_ (.A1(_15478_),
    .A2(_10945_),
    .ZN(_15542_));
 INV_X1 _25257_ (.A(_15542_),
    .ZN(_15543_));
 INV_X1 _25258_ (.A(_15411_),
    .ZN(_15544_));
 AND2_X1 _25259_ (.A1(_15449_),
    .A2(_15410_),
    .ZN(_15545_));
 INV_X2 _25260_ (.A(_15545_),
    .ZN(_15546_));
 OAI22_X1 _25261_ (.A1(_15543_),
    .A2(_15544_),
    .B1(_15546_),
    .B2(_15539_),
    .ZN(_15547_));
 AND2_X1 _25262_ (.A1(_15416_),
    .A2(_10931_),
    .ZN(_15548_));
 AND2_X1 _25263_ (.A1(_15430_),
    .A2(_15548_),
    .ZN(_15549_));
 INV_X1 _25264_ (.A(_15523_),
    .ZN(_15550_));
 AND2_X1 _25265_ (.A1(_15417_),
    .A2(_10945_),
    .ZN(_15551_));
 BUF_X2 _25266_ (.A(_15551_),
    .Z(_15552_));
 INV_X1 _25267_ (.A(_15552_),
    .ZN(_15553_));
 AND2_X2 _25268_ (.A1(_15472_),
    .A2(_10945_),
    .ZN(_15554_));
 INV_X1 _25269_ (.A(_15554_),
    .ZN(_15555_));
 INV_X1 _25270_ (.A(_15498_),
    .ZN(_15556_));
 OAI22_X1 _25271_ (.A1(_15550_),
    .A2(_15553_),
    .B1(_15555_),
    .B2(_15556_),
    .ZN(_15557_));
 NOR4_X1 _25272_ (.A1(_15541_),
    .A2(_15547_),
    .A3(_15549_),
    .A4(_15557_),
    .ZN(_15558_));
 INV_X1 _25273_ (.A(_15415_),
    .ZN(_15559_));
 AND2_X1 _25274_ (.A1(_15505_),
    .A2(_15559_),
    .ZN(_15560_));
 NOR2_X1 _25275_ (.A1(_15455_),
    .A2(_15461_),
    .ZN(_15561_));
 CLKBUF_X2 _25276_ (.A(_15561_),
    .Z(_15562_));
 OAI21_X1 _25277_ (.A(_15532_),
    .B1(_15560_),
    .B2(_15562_),
    .ZN(_15563_));
 AND2_X1 _25278_ (.A1(_15462_),
    .A2(_15415_),
    .ZN(_15564_));
 CLKBUF_X2 _25279_ (.A(_15564_),
    .Z(_15565_));
 INV_X1 _25280_ (.A(_15565_),
    .ZN(_15566_));
 INV_X1 _25281_ (.A(_15497_),
    .ZN(_15567_));
 NAND2_X1 _25282_ (.A1(_15566_),
    .A2(_15567_),
    .ZN(_15568_));
 NOR2_X2 _25283_ (.A1(_15538_),
    .A2(_10964_),
    .ZN(_15569_));
 BUF_X2 _25284_ (.A(_15569_),
    .Z(_15570_));
 NAND2_X1 _25285_ (.A1(_15568_),
    .A2(_15570_),
    .ZN(_15571_));
 CLKBUF_X2 _25286_ (.A(_15491_),
    .Z(_15572_));
 OAI21_X1 _25287_ (.A(_15570_),
    .B1(_15527_),
    .B2(_15572_),
    .ZN(_15573_));
 AND3_X1 _25288_ (.A1(_15563_),
    .A2(_15571_),
    .A3(_15573_),
    .ZN(_15574_));
 AND2_X1 _25289_ (.A1(_15434_),
    .A2(_15532_),
    .ZN(_15575_));
 INV_X1 _25290_ (.A(_15575_),
    .ZN(_15576_));
 AND2_X1 _25291_ (.A1(_15445_),
    .A2(_15440_),
    .ZN(_15577_));
 AND2_X1 _25292_ (.A1(_15478_),
    .A2(_10931_),
    .ZN(_15578_));
 AND2_X1 _25293_ (.A1(_15578_),
    .A2(_15431_),
    .ZN(_15579_));
 NAND2_X1 _25294_ (.A1(_15559_),
    .A2(_15534_),
    .ZN(_15580_));
 NOR2_X1 _25295_ (.A1(_15580_),
    .A2(_15459_),
    .ZN(_15581_));
 AOI211_X1 _25296_ (.A(_15577_),
    .B(_15579_),
    .C1(_15445_),
    .C2(_15581_),
    .ZN(_15582_));
 AND3_X1 _25297_ (.A1(_15574_),
    .A2(_15576_),
    .A3(_15582_),
    .ZN(_15583_));
 NAND4_X1 _25298_ (.A1(_15496_),
    .A2(_15529_),
    .A3(_15558_),
    .A4(_15583_),
    .ZN(_15584_));
 CLKBUF_X2 _25299_ (.A(_15545_),
    .Z(_15585_));
 AND2_X1 _25300_ (.A1(_15462_),
    .A2(_10931_),
    .ZN(_15586_));
 OAI21_X1 _25301_ (.A(_15585_),
    .B1(_15586_),
    .B2(_15520_),
    .ZN(_15587_));
 CLKBUF_X2 _25302_ (.A(_15509_),
    .Z(_15588_));
 AND2_X1 _25303_ (.A1(_15588_),
    .A2(_15520_),
    .ZN(_15589_));
 INV_X1 _25304_ (.A(_15589_),
    .ZN(_15590_));
 AND2_X1 _25305_ (.A1(_15423_),
    .A2(_15462_),
    .ZN(_15591_));
 CLKBUF_X2 _25306_ (.A(_15591_),
    .Z(_15592_));
 OAI21_X1 _25307_ (.A(_15588_),
    .B1(_15592_),
    .B2(_15554_),
    .ZN(_15593_));
 INV_X1 _25308_ (.A(_15534_),
    .ZN(_15594_));
 NOR2_X1 _25309_ (.A1(_15594_),
    .A2(_15486_),
    .ZN(_15595_));
 NAND2_X1 _25310_ (.A1(_15595_),
    .A2(_15513_),
    .ZN(_15596_));
 AND3_X1 _25311_ (.A1(_15590_),
    .A2(_15593_),
    .A3(_15596_),
    .ZN(_15597_));
 BUF_X2 _25312_ (.A(_15417_),
    .Z(_15598_));
 INV_X1 _25313_ (.A(_15475_),
    .ZN(_15599_));
 AND3_X1 _25314_ (.A1(_15585_),
    .A2(_15598_),
    .A3(_15599_),
    .ZN(_15600_));
 OAI21_X1 _25315_ (.A(_15463_),
    .B1(_10932_),
    .B2(_10945_),
    .ZN(_15601_));
 INV_X1 _25316_ (.A(_15601_),
    .ZN(_15602_));
 AOI21_X1 _25317_ (.A(_15600_),
    .B1(_15413_),
    .B2(_15602_),
    .ZN(_15603_));
 CLKBUF_X2 _25318_ (.A(_15507_),
    .Z(_15604_));
 AND2_X1 _25319_ (.A1(_15417_),
    .A2(_15422_),
    .ZN(_15605_));
 OAI21_X1 _25320_ (.A(_15604_),
    .B1(_15586_),
    .B2(_15605_),
    .ZN(_15606_));
 NAND3_X1 _25321_ (.A1(_15507_),
    .A2(_15599_),
    .A3(_15534_),
    .ZN(_15607_));
 AND2_X1 _25322_ (.A1(_15606_),
    .A2(_15607_),
    .ZN(_15608_));
 AND4_X1 _25323_ (.A1(_15587_),
    .A2(_15597_),
    .A3(_15603_),
    .A4(_15608_),
    .ZN(_15609_));
 AND2_X1 _25324_ (.A1(_15506_),
    .A2(_15449_),
    .ZN(_15610_));
 CLKBUF_X2 _25325_ (.A(_15610_),
    .Z(_15611_));
 AND3_X1 _25326_ (.A1(_15611_),
    .A2(_15460_),
    .A3(_15447_),
    .ZN(_15612_));
 AND2_X1 _25327_ (.A1(_15586_),
    .A2(_15471_),
    .ZN(_15613_));
 CLKBUF_X2 _25328_ (.A(_15506_),
    .Z(_15614_));
 AND3_X1 _25329_ (.A1(_15440_),
    .A2(_15614_),
    .A3(_15449_),
    .ZN(_15615_));
 AND2_X1 _25330_ (.A1(_15554_),
    .A2(_15471_),
    .ZN(_15616_));
 NOR4_X1 _25331_ (.A1(_15612_),
    .A2(_15613_),
    .A3(_15615_),
    .A4(_15616_),
    .ZN(_15617_));
 BUF_X2 _25332_ (.A(_15452_),
    .Z(_15618_));
 OAI21_X1 _25333_ (.A(_15618_),
    .B1(_15560_),
    .B2(_15533_),
    .ZN(_15619_));
 AND2_X1 _25334_ (.A1(_15542_),
    .A2(_15484_),
    .ZN(_15620_));
 INV_X1 _25335_ (.A(_15620_),
    .ZN(_15621_));
 AND3_X1 _25336_ (.A1(_15617_),
    .A2(_15619_),
    .A3(_15621_),
    .ZN(_15622_));
 NAND3_X1 _25337_ (.A1(_15505_),
    .A2(_15430_),
    .A3(_15559_),
    .ZN(_15623_));
 NAND2_X1 _25338_ (.A1(_15565_),
    .A2(_15430_),
    .ZN(_15624_));
 AND2_X1 _25339_ (.A1(_15623_),
    .A2(_15624_),
    .ZN(_15625_));
 AND2_X1 _25340_ (.A1(_15474_),
    .A2(_15438_),
    .ZN(_15626_));
 BUF_X2 _25341_ (.A(_15626_),
    .Z(_15627_));
 OAI21_X1 _25342_ (.A(_15522_),
    .B1(_15627_),
    .B2(_15554_),
    .ZN(_15628_));
 NAND4_X1 _25343_ (.A1(_15463_),
    .A2(_15410_),
    .A3(_10932_),
    .A4(_15469_),
    .ZN(_15629_));
 AND2_X1 _25344_ (.A1(_15628_),
    .A2(_15629_),
    .ZN(_15630_));
 INV_X1 _25345_ (.A(_15418_),
    .ZN(_15631_));
 INV_X1 _25346_ (.A(_15433_),
    .ZN(_15632_));
 NAND2_X1 _25347_ (.A1(_15631_),
    .A2(_15632_),
    .ZN(_15633_));
 AND2_X1 _25348_ (.A1(_15438_),
    .A2(_10931_),
    .ZN(_15634_));
 OAI21_X1 _25349_ (.A(_15485_),
    .B1(_15633_),
    .B2(_15634_),
    .ZN(_15635_));
 CLKBUF_X2 _25350_ (.A(_15480_),
    .Z(_15636_));
 BUF_X2 _25351_ (.A(_15636_),
    .Z(_15637_));
 OAI21_X1 _25352_ (.A(_15637_),
    .B1(_15627_),
    .B2(_15533_),
    .ZN(_15638_));
 NAND2_X1 _25353_ (.A1(_15637_),
    .A2(_15456_),
    .ZN(_15639_));
 AND4_X1 _25354_ (.A1(_15630_),
    .A2(_15635_),
    .A3(_15638_),
    .A4(_15639_),
    .ZN(_15640_));
 NAND4_X1 _25355_ (.A1(_15609_),
    .A2(_15622_),
    .A3(_15625_),
    .A4(_15640_),
    .ZN(_15641_));
 NOR2_X2 _25356_ (.A1(_15584_),
    .A2(_15641_),
    .ZN(_15642_));
 XOR2_X1 _25357_ (.A(_15642_),
    .B(_01005_),
    .Z(_15643_));
 MUX2_X1 _25358_ (.A(_01216_),
    .B(_15643_),
    .S(_15147_),
    .Z(_01065_));
 AND2_X1 _25359_ (.A1(_15522_),
    .A2(_15463_),
    .ZN(_15644_));
 AND2_X1 _25360_ (.A1(_15522_),
    .A2(_15627_),
    .ZN(_15645_));
 AND2_X2 _25361_ (.A1(_15424_),
    .A2(_15472_),
    .ZN(_15646_));
 AOI211_X1 _25362_ (.A(_15644_),
    .B(_15645_),
    .C1(_15523_),
    .C2(_15646_),
    .ZN(_15647_));
 INV_X1 _25363_ (.A(_15580_),
    .ZN(_15648_));
 NAND2_X1 _25364_ (.A1(_15648_),
    .A2(_15523_),
    .ZN(_15649_));
 INV_X1 _25365_ (.A(_15548_),
    .ZN(_15650_));
 OAI211_X1 _25366_ (.A(_15647_),
    .B(_15649_),
    .C1(_15650_),
    .C2(_15550_),
    .ZN(_15651_));
 AND2_X1 _25367_ (.A1(_15462_),
    .A2(_10945_),
    .ZN(_15652_));
 AND2_X1 _25368_ (.A1(_15545_),
    .A2(_15652_),
    .ZN(_15653_));
 AND2_X2 _25369_ (.A1(_15478_),
    .A2(_15414_),
    .ZN(_15654_));
 NOR2_X1 _25370_ (.A1(_15654_),
    .A2(_15434_),
    .ZN(_15655_));
 NOR2_X1 _25371_ (.A1(_15655_),
    .A2(_15546_),
    .ZN(_15656_));
 NOR2_X1 _25372_ (.A1(_15520_),
    .A2(_15516_),
    .ZN(_15657_));
 NOR2_X1 _25373_ (.A1(_15657_),
    .A2(_15546_),
    .ZN(_15658_));
 AND2_X1 _25374_ (.A1(_15474_),
    .A2(_15462_),
    .ZN(_15659_));
 AND2_X1 _25375_ (.A1(_15659_),
    .A2(_15545_),
    .ZN(_15660_));
 OR4_X1 _25376_ (.A1(_15653_),
    .A2(_15656_),
    .A3(_15658_),
    .A4(_15660_),
    .ZN(_15661_));
 AND2_X1 _25377_ (.A1(_15411_),
    .A2(_15501_),
    .ZN(_15662_));
 INV_X1 _25378_ (.A(_15662_),
    .ZN(_15663_));
 OAI21_X1 _25379_ (.A(_15412_),
    .B1(_15627_),
    .B2(_15562_),
    .ZN(_15664_));
 AND2_X1 _25380_ (.A1(_15478_),
    .A2(_15422_),
    .ZN(_15665_));
 INV_X1 _25381_ (.A(_15665_),
    .ZN(_15666_));
 OAI211_X1 _25382_ (.A(_15663_),
    .B(_15664_),
    .C1(_15666_),
    .C2(_15544_),
    .ZN(_15667_));
 INV_X1 _25383_ (.A(_15549_),
    .ZN(_15668_));
 NAND4_X1 _25384_ (.A1(_15535_),
    .A2(_15410_),
    .A3(_15429_),
    .A4(_15459_),
    .ZN(_15669_));
 OAI211_X1 _25385_ (.A(_15431_),
    .B(_15464_),
    .C1(_15424_),
    .C2(_15486_),
    .ZN(_15670_));
 NAND2_X1 _25386_ (.A1(_15505_),
    .A2(_15430_),
    .ZN(_15671_));
 NAND4_X1 _25387_ (.A1(_15668_),
    .A2(_15669_),
    .A3(_15670_),
    .A4(_15671_),
    .ZN(_15672_));
 NOR4_X1 _25388_ (.A1(_15651_),
    .A2(_15661_),
    .A3(_15667_),
    .A4(_15672_),
    .ZN(_15673_));
 INV_X1 _25389_ (.A(_15470_),
    .ZN(_15674_));
 INV_X1 _25390_ (.A(_15633_),
    .ZN(_15675_));
 INV_X1 _25391_ (.A(_15578_),
    .ZN(_15676_));
 AOI21_X1 _25392_ (.A(_15674_),
    .B1(_15675_),
    .B2(_15676_),
    .ZN(_15677_));
 AND2_X1 _25393_ (.A1(_15565_),
    .A2(_15471_),
    .ZN(_15678_));
 AND2_X1 _25394_ (.A1(_15516_),
    .A2(_15470_),
    .ZN(_15679_));
 AND2_X1 _25395_ (.A1(_15440_),
    .A2(_15470_),
    .ZN(_15680_));
 NOR4_X1 _25396_ (.A1(_15677_),
    .A2(_15678_),
    .A3(_15679_),
    .A4(_15680_),
    .ZN(_15681_));
 NAND3_X1 _25397_ (.A1(_15516_),
    .A2(_15449_),
    .A3(_15451_),
    .ZN(_15682_));
 INV_X1 _25398_ (.A(_15659_),
    .ZN(_15683_));
 INV_X1 _25399_ (.A(_15453_),
    .ZN(_15684_));
 NAND2_X1 _25400_ (.A1(_15453_),
    .A2(_15439_),
    .ZN(_15685_));
 OAI221_X1 _25401_ (.A(_15682_),
    .B1(_15683_),
    .B2(_15684_),
    .C1(_15436_),
    .C2(_15685_),
    .ZN(_15686_));
 AND4_X1 _25402_ (.A1(_10931_),
    .A2(_15449_),
    .A3(_15417_),
    .A4(_15451_),
    .ZN(_15687_));
 AND2_X1 _25403_ (.A1(_15524_),
    .A2(_15453_),
    .ZN(_15688_));
 NOR4_X1 _25404_ (.A1(_15686_),
    .A2(_15492_),
    .A3(_15687_),
    .A4(_15688_),
    .ZN(_15689_));
 CLKBUF_X2 _25405_ (.A(_15659_),
    .Z(_15690_));
 NAND2_X1 _25406_ (.A1(_15690_),
    .A2(_15484_),
    .ZN(_15691_));
 AND2_X1 _25407_ (.A1(_15483_),
    .A2(_15515_),
    .ZN(_15692_));
 AND3_X1 _25408_ (.A1(_15520_),
    .A2(_15409_),
    .A3(_15451_),
    .ZN(_15693_));
 NOR2_X1 _25409_ (.A1(_15692_),
    .A2(_15693_),
    .ZN(_15694_));
 AND2_X1 _25410_ (.A1(_15652_),
    .A2(_15484_),
    .ZN(_15695_));
 INV_X1 _25411_ (.A(_15695_),
    .ZN(_15696_));
 AND2_X1 _25412_ (.A1(_15526_),
    .A2(_15484_),
    .ZN(_15697_));
 INV_X1 _25413_ (.A(_15697_),
    .ZN(_15698_));
 AND4_X1 _25414_ (.A1(_15691_),
    .A2(_15694_),
    .A3(_15696_),
    .A4(_15698_),
    .ZN(_15699_));
 AND2_X1 _25415_ (.A1(_15565_),
    .A2(_15636_),
    .ZN(_15700_));
 AND2_X1 _25416_ (.A1(_15527_),
    .A2(_15636_),
    .ZN(_15701_));
 AND2_X1 _25417_ (.A1(_15542_),
    .A2(_15636_),
    .ZN(_15702_));
 AND2_X1 _25418_ (.A1(_15636_),
    .A2(_15440_),
    .ZN(_15703_));
 NOR4_X1 _25419_ (.A1(_15700_),
    .A2(_15701_),
    .A3(_15702_),
    .A4(_15703_),
    .ZN(_15704_));
 AND4_X1 _25420_ (.A1(_15681_),
    .A2(_15689_),
    .A3(_15699_),
    .A4(_15704_),
    .ZN(_15705_));
 OAI21_X1 _25421_ (.A(_15531_),
    .B1(_15491_),
    .B2(_15479_),
    .ZN(_15706_));
 NAND3_X1 _25422_ (.A1(_15531_),
    .A2(_15475_),
    .A3(_15534_),
    .ZN(_15707_));
 OAI211_X1 _25423_ (.A(_15706_),
    .B(_15707_),
    .C1(_15537_),
    .C2(_15540_),
    .ZN(_15708_));
 AND3_X1 _25424_ (.A1(_15530_),
    .A2(_15475_),
    .A3(_15463_),
    .ZN(_15709_));
 AND3_X1 _25425_ (.A1(_15530_),
    .A2(_15415_),
    .A3(_15462_),
    .ZN(_15710_));
 OR2_X1 _25426_ (.A1(_15709_),
    .A2(_15710_),
    .ZN(_15711_));
 AND2_X1 _25427_ (.A1(_15554_),
    .A2(_15531_),
    .ZN(_15712_));
 AND2_X1 _25428_ (.A1(_15440_),
    .A2(_15531_),
    .ZN(_15713_));
 NOR4_X1 _25429_ (.A1(_15708_),
    .A2(_15711_),
    .A3(_15712_),
    .A4(_15713_),
    .ZN(_15714_));
 AND2_X1 _25430_ (.A1(_15569_),
    .A2(_15562_),
    .ZN(_15715_));
 INV_X1 _25431_ (.A(_15569_),
    .ZN(_15716_));
 AOI21_X1 _25432_ (.A(_15716_),
    .B1(_15553_),
    .B2(_15666_),
    .ZN(_15717_));
 AOI211_X1 _25433_ (.A(_15715_),
    .B(_15717_),
    .C1(_15570_),
    .C2(_15627_),
    .ZN(_15718_));
 OAI21_X1 _25434_ (.A(_15445_),
    .B1(_15648_),
    .B2(_15514_),
    .ZN(_15719_));
 OAI211_X1 _25435_ (.A(_15498_),
    .B(_15463_),
    .C1(_10931_),
    .C2(_10945_),
    .ZN(_15720_));
 NAND2_X1 _25436_ (.A1(_15626_),
    .A2(_15498_),
    .ZN(_15721_));
 OAI211_X1 _25437_ (.A(_15720_),
    .B(_15721_),
    .C1(_15555_),
    .C2(_15556_),
    .ZN(_15722_));
 AND2_X1 _25438_ (.A1(_15578_),
    .A2(_15498_),
    .ZN(_15723_));
 NOR3_X1 _25439_ (.A1(_15722_),
    .A2(_15502_),
    .A3(_15723_),
    .ZN(_15724_));
 AND4_X1 _25440_ (.A1(_15714_),
    .A2(_15718_),
    .A3(_15719_),
    .A4(_15724_),
    .ZN(_15725_));
 OAI211_X1 _25441_ (.A(_15512_),
    .B(_15472_),
    .C1(_15424_),
    .C2(_15475_),
    .ZN(_15726_));
 OAI21_X1 _25442_ (.A(_15512_),
    .B1(_15527_),
    .B2(_15605_),
    .ZN(_15727_));
 NAND4_X1 _25443_ (.A1(_15614_),
    .A2(_15464_),
    .A3(_10932_),
    .A4(_15429_),
    .ZN(_15728_));
 AND3_X1 _25444_ (.A1(_15726_),
    .A2(_15727_),
    .A3(_15728_),
    .ZN(_15729_));
 AND2_X1 _25445_ (.A1(_15491_),
    .A2(_15509_),
    .ZN(_15730_));
 INV_X1 _25446_ (.A(_15509_),
    .ZN(_15731_));
 INV_X1 _25447_ (.A(_15425_),
    .ZN(_15732_));
 AOI21_X1 _25448_ (.A(_15731_),
    .B1(_15537_),
    .B2(_15732_),
    .ZN(_15733_));
 AOI211_X1 _25449_ (.A(_15730_),
    .B(_15733_),
    .C1(_15602_),
    .C2(_15588_),
    .ZN(_15734_));
 NAND4_X1 _25450_ (.A1(_15614_),
    .A2(_15475_),
    .A3(_15417_),
    .A4(_15469_),
    .ZN(_15735_));
 NAND2_X1 _25451_ (.A1(_15607_),
    .A2(_15735_),
    .ZN(_15736_));
 INV_X1 _25452_ (.A(_15507_),
    .ZN(_15737_));
 INV_X1 _25453_ (.A(_15592_),
    .ZN(_15738_));
 AOI21_X1 _25454_ (.A(_15737_),
    .B1(_15683_),
    .B2(_15738_),
    .ZN(_15739_));
 AOI211_X1 _25455_ (.A(_15736_),
    .B(_15739_),
    .C1(_15520_),
    .C2(_15604_),
    .ZN(_15740_));
 AND2_X1 _25456_ (.A1(_15610_),
    .A2(_15542_),
    .ZN(_15741_));
 AND2_X1 _25457_ (.A1(_15610_),
    .A2(_15493_),
    .ZN(_15742_));
 AND2_X1 _25458_ (.A1(_15610_),
    .A2(_15652_),
    .ZN(_15743_));
 AND2_X1 _25459_ (.A1(_15610_),
    .A2(_15472_),
    .ZN(_15744_));
 NOR4_X1 _25460_ (.A1(_15741_),
    .A2(_15742_),
    .A3(_15743_),
    .A4(_15744_),
    .ZN(_15745_));
 AND4_X1 _25461_ (.A1(_15729_),
    .A2(_15734_),
    .A3(_15740_),
    .A4(_15745_),
    .ZN(_15746_));
 NAND4_X1 _25462_ (.A1(_15673_),
    .A2(_15705_),
    .A3(_15725_),
    .A4(_15746_),
    .ZN(_15747_));
 NOR2_X1 _25463_ (.A1(_15747_),
    .A2(_15575_),
    .ZN(_15748_));
 INV_X1 _25464_ (.A(_01006_),
    .ZN(_15749_));
 XNOR2_X1 _25465_ (.A(_15748_),
    .B(_15749_),
    .ZN(_15750_));
 MUX2_X1 _25466_ (.A(_01217_),
    .B(_15750_),
    .S(_15147_),
    .Z(_01066_));
 AND2_X1 _25467_ (.A1(_15611_),
    .A2(_15565_),
    .ZN(_15751_));
 AND2_X1 _25468_ (.A1(_15611_),
    .A2(_15554_),
    .ZN(_15752_));
 AND2_X1 _25469_ (.A1(_15610_),
    .A2(_15456_),
    .ZN(_15753_));
 NOR4_X1 _25470_ (.A1(_15751_),
    .A2(_15752_),
    .A3(_15753_),
    .A4(_15743_),
    .ZN(_15754_));
 OAI21_X1 _25471_ (.A(_15604_),
    .B1(_15554_),
    .B2(_15533_),
    .ZN(_15755_));
 OAI211_X1 _25472_ (.A(_15604_),
    .B(_15461_),
    .C1(_17068_),
    .C2(_15599_),
    .ZN(_15756_));
 AND3_X1 _25473_ (.A1(_15754_),
    .A2(_15755_),
    .A3(_15756_),
    .ZN(_15757_));
 OAI21_X1 _25474_ (.A(_15512_),
    .B1(_15434_),
    .B2(_15456_),
    .ZN(_15758_));
 AND2_X1 _25475_ (.A1(_15690_),
    .A2(_15588_),
    .ZN(_15759_));
 AOI211_X1 _25476_ (.A(_15594_),
    .B(_15731_),
    .C1(_15437_),
    .C2(_10945_),
    .ZN(_15760_));
 AOI211_X1 _25477_ (.A(_15759_),
    .B(_15760_),
    .C1(_15588_),
    .C2(_15560_),
    .ZN(_15761_));
 AND4_X1 _25478_ (.A1(_15429_),
    .A2(_15614_),
    .A3(_15475_),
    .A4(_15464_),
    .ZN(_15762_));
 INV_X1 _25479_ (.A(_15512_),
    .ZN(_15763_));
 AOI211_X1 _25480_ (.A(_15504_),
    .B(_15763_),
    .C1(_15460_),
    .C2(_15599_),
    .ZN(_15764_));
 AOI211_X1 _25481_ (.A(_15762_),
    .B(_15764_),
    .C1(_15513_),
    .C2(_15652_),
    .ZN(_15765_));
 OAI211_X1 _25482_ (.A(_15513_),
    .B(_15535_),
    .C1(_15437_),
    .C2(_10946_),
    .ZN(_15766_));
 AND4_X1 _25483_ (.A1(_15758_),
    .A2(_15761_),
    .A3(_15765_),
    .A4(_15766_),
    .ZN(_15767_));
 AOI21_X1 _25484_ (.A(_15684_),
    .B1(_15683_),
    .B2(_15738_),
    .ZN(_15768_));
 NAND2_X1 _25485_ (.A1(_15425_),
    .A2(_15453_),
    .ZN(_15769_));
 OAI21_X1 _25486_ (.A(_15769_),
    .B1(_15684_),
    .B2(_15537_),
    .ZN(_15770_));
 NAND2_X1 _25487_ (.A1(_15685_),
    .A2(_15682_),
    .ZN(_15771_));
 OR4_X1 _25488_ (.A1(_15688_),
    .A2(_15768_),
    .A3(_15770_),
    .A4(_15771_),
    .ZN(_15772_));
 AND2_X1 _25489_ (.A1(_15646_),
    .A2(_15471_),
    .ZN(_15773_));
 INV_X1 _25490_ (.A(_15773_),
    .ZN(_15774_));
 OAI211_X1 _25491_ (.A(_15471_),
    .B(_15464_),
    .C1(_10932_),
    .C2(_10938_),
    .ZN(_15775_));
 NAND2_X1 _25492_ (.A1(_15774_),
    .A2(_15775_),
    .ZN(_15776_));
 AND3_X1 _25493_ (.A1(_15535_),
    .A2(_15469_),
    .A3(_15451_),
    .ZN(_15777_));
 AND2_X1 _25494_ (.A1(_15418_),
    .A2(_15470_),
    .ZN(_15778_));
 OR2_X1 _25495_ (.A1(_15494_),
    .A2(_15778_),
    .ZN(_15779_));
 NOR4_X1 _25496_ (.A1(_15772_),
    .A2(_15776_),
    .A3(_15777_),
    .A4(_15779_),
    .ZN(_15780_));
 NAND4_X1 _25497_ (.A1(_15409_),
    .A2(_15473_),
    .A3(_15451_),
    .A4(_10946_),
    .ZN(_15781_));
 OAI21_X1 _25498_ (.A(_15485_),
    .B1(_15690_),
    .B2(_15592_),
    .ZN(_15782_));
 AND2_X1 _25499_ (.A1(_15483_),
    .A2(_15634_),
    .ZN(_15783_));
 INV_X1 _25500_ (.A(_15783_),
    .ZN(_15784_));
 OAI211_X1 _25501_ (.A(_15781_),
    .B(_15782_),
    .C1(_15784_),
    .C2(_10946_),
    .ZN(_15785_));
 INV_X1 _25502_ (.A(_15636_),
    .ZN(_15786_));
 AOI21_X1 _25503_ (.A(_15786_),
    .B1(_15675_),
    .B2(_15543_),
    .ZN(_15787_));
 AND2_X1 _25504_ (.A1(_15524_),
    .A2(_15485_),
    .ZN(_15788_));
 INV_X1 _25505_ (.A(_15561_),
    .ZN(_15789_));
 INV_X1 _25506_ (.A(_15634_),
    .ZN(_15790_));
 AOI21_X1 _25507_ (.A(_15786_),
    .B1(_15789_),
    .B2(_15790_),
    .ZN(_15791_));
 NOR4_X1 _25508_ (.A1(_15785_),
    .A2(_15787_),
    .A3(_15788_),
    .A4(_15791_),
    .ZN(_15792_));
 AND4_X1 _25509_ (.A1(_15757_),
    .A2(_15767_),
    .A3(_15780_),
    .A4(_15792_),
    .ZN(_15793_));
 OAI211_X1 _25510_ (.A(_15570_),
    .B(_15533_),
    .C1(_10932_),
    .C2(_10946_),
    .ZN(_15794_));
 OAI21_X1 _25511_ (.A(_15570_),
    .B1(_15527_),
    .B2(_15419_),
    .ZN(_15795_));
 OAI211_X1 _25512_ (.A(_15794_),
    .B(_15795_),
    .C1(_15555_),
    .C2(_15716_),
    .ZN(_15796_));
 NOR2_X1 _25513_ (.A1(_15504_),
    .A2(_15474_),
    .ZN(_15797_));
 NAND2_X1 _25514_ (.A1(_15797_),
    .A2(_15530_),
    .ZN(_15798_));
 NAND3_X1 _25515_ (.A1(_15530_),
    .A2(_15475_),
    .A3(_15463_),
    .ZN(_15799_));
 NAND2_X1 _25516_ (.A1(_15798_),
    .A2(_15799_),
    .ZN(_15800_));
 AND2_X1 _25517_ (.A1(_15524_),
    .A2(_15532_),
    .ZN(_15801_));
 AND3_X1 _25518_ (.A1(_15501_),
    .A2(_15559_),
    .A3(_15532_),
    .ZN(_15802_));
 NOR4_X1 _25519_ (.A1(_15796_),
    .A2(_15800_),
    .A3(_15801_),
    .A4(_15802_),
    .ZN(_15803_));
 OAI21_X1 _25520_ (.A(_15413_),
    .B1(_15568_),
    .B2(_15560_),
    .ZN(_15804_));
 AND2_X1 _25521_ (.A1(_15431_),
    .A2(_15646_),
    .ZN(_15805_));
 AND2_X1 _25522_ (.A1(_15652_),
    .A2(_15430_),
    .ZN(_15806_));
 AND2_X1 _25523_ (.A1(_15431_),
    .A2(_15419_),
    .ZN(_15807_));
 NOR4_X1 _25524_ (.A1(_15579_),
    .A2(_15805_),
    .A3(_15806_),
    .A4(_15807_),
    .ZN(_15808_));
 OAI21_X1 _25525_ (.A(_15523_),
    .B1(_15572_),
    .B2(_15493_),
    .ZN(_15809_));
 OAI21_X1 _25526_ (.A(_15523_),
    .B1(_15690_),
    .B2(_15440_),
    .ZN(_15810_));
 OAI21_X1 _25527_ (.A(_15585_),
    .B1(_15572_),
    .B2(_15419_),
    .ZN(_15811_));
 OAI21_X1 _25528_ (.A(_15585_),
    .B1(_15690_),
    .B2(_15634_),
    .ZN(_15812_));
 AND4_X1 _25529_ (.A1(_15809_),
    .A2(_15810_),
    .A3(_15811_),
    .A4(_15812_),
    .ZN(_15813_));
 AND2_X1 _25530_ (.A1(_15413_),
    .A2(_15654_),
    .ZN(_15814_));
 AND2_X1 _25531_ (.A1(_15572_),
    .A2(_15412_),
    .ZN(_15815_));
 NOR3_X1 _25532_ (.A1(_15814_),
    .A2(_15815_),
    .A3(_15426_),
    .ZN(_15816_));
 AND4_X1 _25533_ (.A1(_15804_),
    .A2(_15808_),
    .A3(_15813_),
    .A4(_15816_),
    .ZN(_15817_));
 NAND4_X1 _25534_ (.A1(_15486_),
    .A2(_15409_),
    .A3(_15464_),
    .A4(_15443_),
    .ZN(_15818_));
 NAND4_X1 _25535_ (.A1(_15409_),
    .A2(_15473_),
    .A3(_15415_),
    .A4(_15443_),
    .ZN(_15819_));
 INV_X1 _25536_ (.A(_15444_),
    .ZN(_15820_));
 INV_X1 _25537_ (.A(_15652_),
    .ZN(_15821_));
 OAI211_X1 _25538_ (.A(_15818_),
    .B(_15819_),
    .C1(_15820_),
    .C2(_15821_),
    .ZN(_15822_));
 NAND2_X1 _25539_ (.A1(_15599_),
    .A2(_15598_),
    .ZN(_15823_));
 NOR2_X1 _25540_ (.A1(_15820_),
    .A2(_15823_),
    .ZN(_15824_));
 AND2_X1 _25541_ (.A1(_15445_),
    .A2(_15542_),
    .ZN(_15825_));
 AND2_X1 _25542_ (.A1(_15445_),
    .A2(_15524_),
    .ZN(_15826_));
 NOR4_X1 _25543_ (.A1(_15822_),
    .A2(_15824_),
    .A3(_15825_),
    .A4(_15826_),
    .ZN(_15827_));
 OAI21_X1 _25544_ (.A(_15499_),
    .B1(_15581_),
    .B2(_15552_),
    .ZN(_15828_));
 OAI21_X1 _25545_ (.A(_15499_),
    .B1(_15497_),
    .B2(_15634_),
    .ZN(_15829_));
 AND2_X1 _25546_ (.A1(_15828_),
    .A2(_15829_),
    .ZN(_15830_));
 AND4_X1 _25547_ (.A1(_15803_),
    .A2(_15817_),
    .A3(_15827_),
    .A4(_15830_),
    .ZN(_15831_));
 AND2_X1 _25548_ (.A1(_15793_),
    .A2(_15831_),
    .ZN(_15832_));
 XOR2_X1 _25549_ (.A(_15832_),
    .B(_01007_),
    .Z(_15833_));
 MUX2_X1 _25550_ (.A(_01218_),
    .B(_15833_),
    .S(_15147_),
    .Z(_01067_));
 OAI21_X1 _25551_ (.A(_15532_),
    .B1(_15581_),
    .B2(_15548_),
    .ZN(_15834_));
 AND2_X1 _25552_ (.A1(_15627_),
    .A2(_15531_),
    .ZN(_15835_));
 AND2_X1 _25553_ (.A1(_15516_),
    .A2(_15532_),
    .ZN(_15836_));
 NOR3_X1 _25554_ (.A1(_15835_),
    .A2(_15710_),
    .A3(_15836_),
    .ZN(_15837_));
 OAI21_X1 _25555_ (.A(_15570_),
    .B1(_15568_),
    .B2(_15516_),
    .ZN(_15838_));
 OAI21_X1 _25556_ (.A(_15570_),
    .B1(_15493_),
    .B2(_15419_),
    .ZN(_15839_));
 NAND2_X1 _25557_ (.A1(_15542_),
    .A2(_15569_),
    .ZN(_15840_));
 NAND4_X1 _25558_ (.A1(_15449_),
    .A2(_15459_),
    .A3(_15598_),
    .A4(_15443_),
    .ZN(_15841_));
 AND3_X1 _25559_ (.A1(_15839_),
    .A2(_15840_),
    .A3(_15841_),
    .ZN(_15842_));
 AND4_X1 _25560_ (.A1(_15834_),
    .A2(_15837_),
    .A3(_15838_),
    .A4(_15842_),
    .ZN(_15843_));
 AOI211_X1 _25561_ (.A(_15504_),
    .B(_15544_),
    .C1(_15437_),
    .C2(_10946_),
    .ZN(_15844_));
 AND2_X1 _25562_ (.A1(_15412_),
    .A2(_15586_),
    .ZN(_15845_));
 OR4_X1 _25563_ (.A1(_15662_),
    .A2(_15844_),
    .A3(_15815_),
    .A4(_15845_),
    .ZN(_15846_));
 AND4_X1 _25564_ (.A1(_15460_),
    .A2(_15431_),
    .A3(_15559_),
    .A4(_15535_),
    .ZN(_15847_));
 INV_X1 _25565_ (.A(_15430_),
    .ZN(_15848_));
 AND2_X1 _25566_ (.A1(_15463_),
    .A2(_15422_),
    .ZN(_15849_));
 INV_X1 _25567_ (.A(_15849_),
    .ZN(_15850_));
 INV_X1 _25568_ (.A(_15646_),
    .ZN(_15851_));
 AOI21_X1 _25569_ (.A(_15848_),
    .B1(_15850_),
    .B2(_15851_),
    .ZN(_15852_));
 NOR4_X1 _25570_ (.A1(_15846_),
    .A2(_15807_),
    .A3(_15847_),
    .A4(_15852_),
    .ZN(_15853_));
 OR2_X1 _25571_ (.A1(_15479_),
    .A2(_15654_),
    .ZN(_15854_));
 AND2_X1 _25572_ (.A1(_15854_),
    .A2(_15499_),
    .ZN(_15855_));
 AND2_X1 _25573_ (.A1(_15515_),
    .A2(_15498_),
    .ZN(_15856_));
 AOI21_X1 _25574_ (.A(_15820_),
    .B1(_15732_),
    .B2(_15676_),
    .ZN(_15857_));
 AND2_X1 _25575_ (.A1(_15444_),
    .A2(_15646_),
    .ZN(_15858_));
 NOR4_X1 _25576_ (.A1(_15855_),
    .A2(_15856_),
    .A3(_15857_),
    .A4(_15858_),
    .ZN(_15859_));
 AOI21_X1 _25577_ (.A(_15546_),
    .B1(_15631_),
    .B2(_15676_),
    .ZN(_15860_));
 AND2_X1 _25578_ (.A1(_15585_),
    .A2(_15562_),
    .ZN(_15861_));
 AND2_X1 _25579_ (.A1(_15545_),
    .A2(_15472_),
    .ZN(_15862_));
 NOR4_X1 _25580_ (.A1(_15860_),
    .A2(_15653_),
    .A3(_15861_),
    .A4(_15862_),
    .ZN(_15863_));
 OAI211_X1 _25581_ (.A(_15523_),
    .B(_15598_),
    .C1(_15437_),
    .C2(_10938_),
    .ZN(_15864_));
 AND2_X1 _25582_ (.A1(_15472_),
    .A2(_15422_),
    .ZN(_15865_));
 OAI21_X1 _25583_ (.A(_15523_),
    .B1(_15592_),
    .B2(_15865_),
    .ZN(_15866_));
 AND4_X1 _25584_ (.A1(_15649_),
    .A2(_15863_),
    .A3(_15864_),
    .A4(_15866_),
    .ZN(_15867_));
 AND4_X1 _25585_ (.A1(_15843_),
    .A2(_15853_),
    .A3(_15859_),
    .A4(_15867_),
    .ZN(_15868_));
 AND4_X1 _25586_ (.A1(_10938_),
    .A2(_15614_),
    .A3(_15429_),
    .A4(_15473_),
    .ZN(_15869_));
 AND2_X1 _25587_ (.A1(_15512_),
    .A2(_15646_),
    .ZN(_15870_));
 AOI211_X1 _25588_ (.A(_15869_),
    .B(_15870_),
    .C1(_15513_),
    .C2(_15568_),
    .ZN(_15871_));
 NAND4_X1 _25589_ (.A1(_15614_),
    .A2(_10932_),
    .A3(_15429_),
    .A4(_15598_),
    .ZN(_15872_));
 OAI211_X1 _25590_ (.A(_15513_),
    .B(_15535_),
    .C1(_15437_),
    .C2(_10938_),
    .ZN(_15873_));
 AND3_X1 _25591_ (.A1(_15871_),
    .A2(_15872_),
    .A3(_15873_),
    .ZN(_15874_));
 NOR2_X1 _25592_ (.A1(_15737_),
    .A2(_15823_),
    .ZN(_15875_));
 AND3_X1 _25593_ (.A1(_15505_),
    .A2(_15604_),
    .A3(_15559_),
    .ZN(_15876_));
 AND2_X1 _25594_ (.A1(_15479_),
    .A2(_15604_),
    .ZN(_15877_));
 AND2_X1 _25595_ (.A1(_15604_),
    .A2(_15562_),
    .ZN(_15878_));
 NOR4_X1 _25596_ (.A1(_15875_),
    .A2(_15876_),
    .A3(_15877_),
    .A4(_15878_),
    .ZN(_15879_));
 NOR2_X1 _25597_ (.A1(_15690_),
    .A2(_15591_),
    .ZN(_15880_));
 INV_X1 _25598_ (.A(_15610_),
    .ZN(_15881_));
 NOR2_X1 _25599_ (.A1(_15880_),
    .A2(_15881_),
    .ZN(_15882_));
 AND2_X1 _25600_ (.A1(_15611_),
    .A2(_15578_),
    .ZN(_15883_));
 NOR4_X1 _25601_ (.A1(_15882_),
    .A2(_15744_),
    .A3(_15753_),
    .A4(_15883_),
    .ZN(_15884_));
 AND2_X1 _25602_ (.A1(_15509_),
    .A2(_15654_),
    .ZN(_15885_));
 NOR2_X1 _25603_ (.A1(_15510_),
    .A2(_15885_),
    .ZN(_15886_));
 INV_X1 _25604_ (.A(_15886_),
    .ZN(_15887_));
 AND2_X1 _25605_ (.A1(_15588_),
    .A2(_15456_),
    .ZN(_15888_));
 NOR4_X1 _25606_ (.A1(_15887_),
    .A2(_15589_),
    .A3(_15888_),
    .A4(_15759_),
    .ZN(_15889_));
 NAND4_X1 _25607_ (.A1(_15874_),
    .A2(_15879_),
    .A3(_15884_),
    .A4(_15889_),
    .ZN(_15890_));
 INV_X1 _25608_ (.A(_15778_),
    .ZN(_15891_));
 NAND3_X1 _25609_ (.A1(_15471_),
    .A2(_15459_),
    .A3(_15535_),
    .ZN(_15892_));
 OAI211_X1 _25610_ (.A(_15891_),
    .B(_15892_),
    .C1(_15553_),
    .C2(_15674_),
    .ZN(_15893_));
 AOI21_X1 _25611_ (.A(_15674_),
    .B1(_15566_),
    .B2(_15821_),
    .ZN(_15894_));
 NOR4_X1 _25612_ (.A1(_15893_),
    .A2(_15616_),
    .A3(_15680_),
    .A4(_15894_),
    .ZN(_15895_));
 NAND2_X1 _25613_ (.A1(_15565_),
    .A2(_15453_),
    .ZN(_15896_));
 OAI21_X1 _25614_ (.A(_15618_),
    .B1(_15479_),
    .B2(_15654_),
    .ZN(_15897_));
 AND4_X1 _25615_ (.A1(_15896_),
    .A2(_15897_),
    .A3(_15685_),
    .A4(_15769_),
    .ZN(_15898_));
 NAND2_X1 _25616_ (.A1(_15895_),
    .A2(_15898_),
    .ZN(_15899_));
 OAI211_X1 _25617_ (.A(_15485_),
    .B(_15598_),
    .C1(_15424_),
    .C2(_15486_),
    .ZN(_15900_));
 OAI211_X1 _25618_ (.A(_15485_),
    .B(_15535_),
    .C1(_15437_),
    .C2(_10946_),
    .ZN(_15901_));
 OAI211_X1 _25619_ (.A(_15485_),
    .B(_15533_),
    .C1(_10932_),
    .C2(_10946_),
    .ZN(_15902_));
 OAI21_X1 _25620_ (.A(_15485_),
    .B1(_15516_),
    .B2(_15440_),
    .ZN(_15903_));
 NAND4_X1 _25621_ (.A1(_15900_),
    .A2(_15901_),
    .A3(_15902_),
    .A4(_15903_),
    .ZN(_15904_));
 OAI211_X1 _25622_ (.A(_15637_),
    .B(_15535_),
    .C1(_15459_),
    .C2(_15415_),
    .ZN(_15905_));
 OAI211_X1 _25623_ (.A(_15637_),
    .B(_15533_),
    .C1(_10938_),
    .C2(_15424_),
    .ZN(_15906_));
 NAND3_X1 _25624_ (.A1(_15637_),
    .A2(_15473_),
    .A3(_15486_),
    .ZN(_15907_));
 OAI21_X1 _25625_ (.A(_15637_),
    .B1(_15434_),
    .B2(_15456_),
    .ZN(_15908_));
 NAND4_X1 _25626_ (.A1(_15905_),
    .A2(_15906_),
    .A3(_15907_),
    .A4(_15908_),
    .ZN(_15909_));
 NOR4_X1 _25627_ (.A1(_15890_),
    .A2(_15899_),
    .A3(_15904_),
    .A4(_15909_),
    .ZN(_15910_));
 AND2_X1 _25628_ (.A1(_15868_),
    .A2(_15910_),
    .ZN(_15911_));
 INV_X1 _25629_ (.A(_01008_),
    .ZN(_15912_));
 XNOR2_X1 _25630_ (.A(_15911_),
    .B(_15912_),
    .ZN(_15913_));
 MUX2_X1 _25631_ (.A(_01219_),
    .B(_15913_),
    .S(_15147_),
    .Z(_01068_));
 NAND3_X1 _25632_ (.A1(_15532_),
    .A2(_15459_),
    .A3(_15533_),
    .ZN(_15914_));
 AOI211_X1 _25633_ (.A(_15504_),
    .B(_15716_),
    .C1(_15460_),
    .C2(_15599_),
    .ZN(_15915_));
 AND2_X1 _25634_ (.A1(_15569_),
    .A2(_15418_),
    .ZN(_15916_));
 AND2_X1 _25635_ (.A1(_15592_),
    .A2(_15569_),
    .ZN(_15917_));
 INV_X1 _25636_ (.A(_15654_),
    .ZN(_15918_));
 OAI21_X1 _25637_ (.A(_15840_),
    .B1(_15918_),
    .B2(_15716_),
    .ZN(_15919_));
 NOR4_X1 _25638_ (.A1(_15915_),
    .A2(_15916_),
    .A3(_15917_),
    .A4(_15919_),
    .ZN(_15920_));
 OAI21_X1 _25639_ (.A(_15532_),
    .B1(_15479_),
    .B2(_15501_),
    .ZN(_15921_));
 AND4_X1 _25640_ (.A1(_15914_),
    .A2(_15920_),
    .A3(_15798_),
    .A4(_15921_),
    .ZN(_15922_));
 NAND2_X1 _25641_ (.A1(_15595_),
    .A2(_15499_),
    .ZN(_15923_));
 AND2_X1 _25642_ (.A1(_15444_),
    .A2(_15554_),
    .ZN(_15924_));
 AOI211_X1 _25643_ (.A(_15577_),
    .B(_15924_),
    .C1(_15445_),
    .C2(_15568_),
    .ZN(_15925_));
 OAI21_X1 _25644_ (.A(_15445_),
    .B1(_15648_),
    .B2(_15447_),
    .ZN(_15926_));
 INV_X1 _25645_ (.A(_15520_),
    .ZN(_15927_));
 OAI21_X1 _25646_ (.A(_15721_),
    .B1(_15927_),
    .B2(_15556_),
    .ZN(_15928_));
 AND2_X1 _25647_ (.A1(_15592_),
    .A2(_15499_),
    .ZN(_15929_));
 NOR2_X1 _25648_ (.A1(_15928_),
    .A2(_15929_),
    .ZN(_15930_));
 AND4_X1 _25649_ (.A1(_15923_),
    .A2(_15925_),
    .A3(_15926_),
    .A4(_15930_),
    .ZN(_15931_));
 NAND2_X1 _25650_ (.A1(_15572_),
    .A2(_15585_),
    .ZN(_15932_));
 NAND2_X1 _25651_ (.A1(_15585_),
    .A2(_15552_),
    .ZN(_15933_));
 OAI211_X1 _25652_ (.A(_15932_),
    .B(_15933_),
    .C1(_15539_),
    .C2(_15546_),
    .ZN(_15934_));
 AOI21_X1 _25653_ (.A(_15550_),
    .B1(_15631_),
    .B2(_15666_),
    .ZN(_15935_));
 NAND2_X1 _25654_ (.A1(_15585_),
    .A2(_15627_),
    .ZN(_15936_));
 OAI21_X1 _25655_ (.A(_15936_),
    .B1(_15546_),
    .B2(_15789_),
    .ZN(_15937_));
 NOR4_X1 _25656_ (.A1(_15934_),
    .A2(_15935_),
    .A3(_15937_),
    .A4(_15644_),
    .ZN(_15938_));
 INV_X1 _25657_ (.A(_15845_),
    .ZN(_15939_));
 NAND2_X1 _25658_ (.A1(_15527_),
    .A2(_15412_),
    .ZN(_15940_));
 OAI21_X1 _25659_ (.A(_15413_),
    .B1(_15419_),
    .B2(_15434_),
    .ZN(_15941_));
 OAI211_X1 _25660_ (.A(_15413_),
    .B(_15473_),
    .C1(_15437_),
    .C2(_10946_),
    .ZN(_15942_));
 NAND4_X1 _25661_ (.A1(_15939_),
    .A2(_15940_),
    .A3(_15941_),
    .A4(_15942_),
    .ZN(_15943_));
 AND2_X1 _25662_ (.A1(_15690_),
    .A2(_15431_),
    .ZN(_15944_));
 OR2_X1 _25663_ (.A1(_15806_),
    .A2(_15944_),
    .ZN(_15945_));
 AND2_X1 _25664_ (.A1(_15431_),
    .A2(_15473_),
    .ZN(_15946_));
 NAND2_X1 _25665_ (.A1(_15542_),
    .A2(_15431_),
    .ZN(_15947_));
 OAI211_X1 _25666_ (.A(_15947_),
    .B(_15435_),
    .C1(_15539_),
    .C2(_15848_),
    .ZN(_15948_));
 NOR4_X1 _25667_ (.A1(_15943_),
    .A2(_15945_),
    .A3(_15946_),
    .A4(_15948_),
    .ZN(_15949_));
 NAND4_X1 _25668_ (.A1(_15922_),
    .A2(_15931_),
    .A3(_15938_),
    .A4(_15949_),
    .ZN(_15950_));
 AND2_X1 _25669_ (.A1(_15592_),
    .A2(_15636_),
    .ZN(_15951_));
 AOI211_X1 _25670_ (.A(_15481_),
    .B(_15951_),
    .C1(_15473_),
    .C2(_15637_),
    .ZN(_15952_));
 OAI21_X1 _25671_ (.A(_15485_),
    .B1(_15578_),
    .B2(_15501_),
    .ZN(_15953_));
 AND4_X1 _25672_ (.A1(_15784_),
    .A2(_15952_),
    .A3(_15696_),
    .A4(_15953_),
    .ZN(_15954_));
 INV_X1 _25673_ (.A(_15870_),
    .ZN(_15955_));
 INV_X1 _25674_ (.A(_15885_),
    .ZN(_15956_));
 OAI211_X1 _25675_ (.A(_15588_),
    .B(_15598_),
    .C1(_15424_),
    .C2(_15486_),
    .ZN(_15957_));
 AND4_X1 _25676_ (.A1(_15590_),
    .A2(_15956_),
    .A3(_15593_),
    .A4(_15957_),
    .ZN(_15958_));
 OAI21_X1 _25677_ (.A(_15513_),
    .B1(_15690_),
    .B2(_15592_),
    .ZN(_15959_));
 OAI21_X1 _25678_ (.A(_15513_),
    .B1(_15572_),
    .B2(_15493_),
    .ZN(_15960_));
 AND4_X1 _25679_ (.A1(_15955_),
    .A2(_15958_),
    .A3(_15959_),
    .A4(_15960_),
    .ZN(_15961_));
 OAI21_X1 _25680_ (.A(_15611_),
    .B1(_15527_),
    .B2(_15419_),
    .ZN(_15962_));
 NAND4_X1 _25681_ (.A1(_15614_),
    .A2(_15533_),
    .A3(_15449_),
    .A4(_10938_),
    .ZN(_15963_));
 NAND2_X1 _25682_ (.A1(_15797_),
    .A2(_15611_),
    .ZN(_15964_));
 NAND3_X1 _25683_ (.A1(_15962_),
    .A2(_15963_),
    .A3(_15964_),
    .ZN(_15965_));
 NOR4_X1 _25684_ (.A1(_15965_),
    .A2(_15736_),
    .A3(_15508_),
    .A4(_15878_),
    .ZN(_15966_));
 OAI21_X1 _25685_ (.A(_15618_),
    .B1(_15592_),
    .B2(_15562_),
    .ZN(_15967_));
 OAI21_X1 _25686_ (.A(_15618_),
    .B1(_15493_),
    .B2(_15552_),
    .ZN(_15968_));
 NAND2_X1 _25687_ (.A1(_15527_),
    .A2(_15618_),
    .ZN(_15969_));
 NAND4_X1 _25688_ (.A1(_15967_),
    .A2(_15968_),
    .A3(_15685_),
    .A4(_15969_),
    .ZN(_15970_));
 AOI21_X1 _25689_ (.A(_15674_),
    .B1(_15666_),
    .B2(_15553_),
    .ZN(_15971_));
 NOR3_X1 _25690_ (.A1(_15776_),
    .A2(_15970_),
    .A3(_15971_),
    .ZN(_15972_));
 NAND4_X1 _25691_ (.A1(_15954_),
    .A2(_15961_),
    .A3(_15966_),
    .A4(_15972_),
    .ZN(_15973_));
 NOR2_X1 _25692_ (.A1(_15950_),
    .A2(_15973_),
    .ZN(_15974_));
 XOR2_X1 _25693_ (.A(_15974_),
    .B(_01009_),
    .Z(_15975_));
 MUX2_X1 _25694_ (.A(_01220_),
    .B(_15975_),
    .S(_15147_),
    .Z(_01070_));
 AND4_X1 _25695_ (.A1(_15460_),
    .A2(_15470_),
    .A3(_15559_),
    .A4(_15534_),
    .ZN(_15976_));
 AOI211_X1 _25696_ (.A(_15976_),
    .B(_15779_),
    .C1(_15552_),
    .C2(_15471_),
    .ZN(_15977_));
 OAI21_X1 _25697_ (.A(_15484_),
    .B1(_15627_),
    .B2(_15565_),
    .ZN(_15978_));
 NAND2_X1 _25698_ (.A1(_15491_),
    .A2(_15636_),
    .ZN(_15979_));
 NAND2_X1 _25699_ (.A1(_15654_),
    .A2(_15636_),
    .ZN(_15980_));
 AND4_X1 _25700_ (.A1(_15482_),
    .A2(_15979_),
    .A3(_15489_),
    .A4(_15980_),
    .ZN(_15981_));
 OAI21_X1 _25701_ (.A(_15484_),
    .B1(_15479_),
    .B2(_15552_),
    .ZN(_15982_));
 OAI21_X1 _25702_ (.A(_15636_),
    .B1(_15690_),
    .B2(_15865_),
    .ZN(_15983_));
 AND4_X1 _25703_ (.A1(_15978_),
    .A2(_15981_),
    .A3(_15982_),
    .A4(_15983_),
    .ZN(_15984_));
 OAI21_X1 _25704_ (.A(_15471_),
    .B1(_15849_),
    .B2(_15646_),
    .ZN(_15985_));
 OAI21_X1 _25705_ (.A(_15896_),
    .B1(_15821_),
    .B2(_15684_),
    .ZN(_15986_));
 AND2_X1 _25706_ (.A1(_15526_),
    .A2(_15453_),
    .ZN(_15987_));
 AND2_X1 _25707_ (.A1(_15453_),
    .A2(_15552_),
    .ZN(_15988_));
 NOR4_X1 _25708_ (.A1(_15986_),
    .A2(_15457_),
    .A3(_15987_),
    .A4(_15988_),
    .ZN(_15989_));
 AND4_X1 _25709_ (.A1(_15977_),
    .A2(_15984_),
    .A3(_15985_),
    .A4(_15989_),
    .ZN(_15990_));
 AND2_X1 _25710_ (.A1(_15554_),
    .A2(_15498_),
    .ZN(_15991_));
 NOR2_X1 _25711_ (.A1(_15928_),
    .A2(_15991_),
    .ZN(_15992_));
 NAND2_X1 _25712_ (.A1(_15565_),
    .A2(_15499_),
    .ZN(_15993_));
 NAND4_X1 _25713_ (.A1(_15486_),
    .A2(_15429_),
    .A3(_15598_),
    .A4(_15443_),
    .ZN(_15994_));
 AND3_X1 _25714_ (.A1(_15992_),
    .A2(_15993_),
    .A3(_15994_),
    .ZN(_15995_));
 NAND2_X1 _25715_ (.A1(_15444_),
    .A2(_15562_),
    .ZN(_15996_));
 NAND4_X1 _25716_ (.A1(_15409_),
    .A2(_15436_),
    .A3(_15472_),
    .A4(_15443_),
    .ZN(_15997_));
 OAI211_X1 _25717_ (.A(_15996_),
    .B(_15997_),
    .C1(_15820_),
    .C2(_15821_),
    .ZN(_15998_));
 AOI211_X1 _25718_ (.A(_15824_),
    .B(_15998_),
    .C1(_15445_),
    .C2(_15648_),
    .ZN(_15999_));
 AND2_X1 _25719_ (.A1(_15854_),
    .A2(_15569_),
    .ZN(_16000_));
 AND3_X1 _25720_ (.A1(_15505_),
    .A2(_15569_),
    .A3(_15559_),
    .ZN(_16001_));
 AOI21_X1 _25721_ (.A(_15716_),
    .B1(_15789_),
    .B2(_15567_),
    .ZN(_16002_));
 NOR4_X1 _25722_ (.A1(_16000_),
    .A2(_15916_),
    .A3(_16001_),
    .A4(_16002_),
    .ZN(_16003_));
 NAND2_X1 _25723_ (.A1(_15501_),
    .A2(_15531_),
    .ZN(_16004_));
 OAI221_X1 _25724_ (.A(_15531_),
    .B1(_15436_),
    .B2(_10938_),
    .C1(_15472_),
    .C2(_15463_),
    .ZN(_16005_));
 AND4_X1 _25725_ (.A1(_16004_),
    .A2(_15706_),
    .A3(_16005_),
    .A4(_15707_),
    .ZN(_16006_));
 AND4_X1 _25726_ (.A1(_15995_),
    .A2(_15999_),
    .A3(_16003_),
    .A4(_16006_),
    .ZN(_16007_));
 AOI21_X1 _25727_ (.A(_15546_),
    .B1(_15789_),
    .B2(_15567_),
    .ZN(_16008_));
 NAND2_X1 _25728_ (.A1(_15527_),
    .A2(_15585_),
    .ZN(_16009_));
 OAI21_X1 _25729_ (.A(_16009_),
    .B1(_15546_),
    .B2(_15543_),
    .ZN(_16010_));
 AND2_X1 _25730_ (.A1(_15585_),
    .A2(_15419_),
    .ZN(_16011_));
 NOR3_X1 _25731_ (.A1(_16008_),
    .A2(_16010_),
    .A3(_16011_),
    .ZN(_16012_));
 NAND2_X1 _25732_ (.A1(_15412_),
    .A2(_15634_),
    .ZN(_16013_));
 AND4_X1 _25733_ (.A1(_15940_),
    .A2(_15939_),
    .A3(_15663_),
    .A4(_16013_),
    .ZN(_16014_));
 INV_X1 _25734_ (.A(_15806_),
    .ZN(_16015_));
 OAI21_X1 _25735_ (.A(_15430_),
    .B1(_15425_),
    .B2(_15524_),
    .ZN(_16016_));
 AND4_X1 _25736_ (.A1(_15624_),
    .A2(_16015_),
    .A3(_15623_),
    .A4(_16016_),
    .ZN(_16017_));
 OAI21_X1 _25737_ (.A(_15522_),
    .B1(_15493_),
    .B2(_15578_),
    .ZN(_16018_));
 AND3_X1 _25738_ (.A1(_16018_),
    .A2(_15629_),
    .A3(_15628_),
    .ZN(_16019_));
 AND4_X1 _25739_ (.A1(_16012_),
    .A2(_16014_),
    .A3(_16017_),
    .A4(_16019_),
    .ZN(_16020_));
 AND2_X1 _25740_ (.A1(_15507_),
    .A2(_15419_),
    .ZN(_16021_));
 AOI21_X1 _25741_ (.A(_15737_),
    .B1(_15738_),
    .B2(_15789_),
    .ZN(_16022_));
 INV_X1 _25742_ (.A(_15657_),
    .ZN(_16023_));
 AOI211_X1 _25743_ (.A(_16021_),
    .B(_16022_),
    .C1(_15604_),
    .C2(_16023_),
    .ZN(_16024_));
 AOI211_X1 _25744_ (.A(_15741_),
    .B(_15882_),
    .C1(_15434_),
    .C2(_15611_),
    .ZN(_16025_));
 AOI21_X1 _25745_ (.A(_15731_),
    .B1(_15683_),
    .B2(_15566_),
    .ZN(_16026_));
 OAI211_X1 _25746_ (.A(_15509_),
    .B(_15598_),
    .C1(_15436_),
    .C2(_10945_),
    .ZN(_16027_));
 INV_X1 _25747_ (.A(_16027_),
    .ZN(_16028_));
 AND2_X1 _25748_ (.A1(_15509_),
    .A2(_15440_),
    .ZN(_16029_));
 AND2_X1 _25749_ (.A1(_15526_),
    .A2(_15509_),
    .ZN(_16030_));
 NOR4_X1 _25750_ (.A1(_16026_),
    .A2(_16028_),
    .A3(_16029_),
    .A4(_16030_),
    .ZN(_16031_));
 NAND2_X1 _25751_ (.A1(_15512_),
    .A2(_15654_),
    .ZN(_16032_));
 OAI211_X1 _25752_ (.A(_15511_),
    .B(_15472_),
    .C1(_15436_),
    .C2(_10945_),
    .ZN(_16033_));
 OAI21_X1 _25753_ (.A(_15512_),
    .B1(_15497_),
    .B2(_15562_),
    .ZN(_16034_));
 AND4_X1 _25754_ (.A1(_16032_),
    .A2(_16033_),
    .A3(_15758_),
    .A4(_16034_),
    .ZN(_16035_));
 AND4_X1 _25755_ (.A1(_16024_),
    .A2(_16025_),
    .A3(_16031_),
    .A4(_16035_),
    .ZN(_16036_));
 NAND4_X1 _25756_ (.A1(_15990_),
    .A2(_16007_),
    .A3(_16020_),
    .A4(_16036_),
    .ZN(_16037_));
 NOR2_X1 _25757_ (.A1(_16037_),
    .A2(_15575_),
    .ZN(_16038_));
 XOR2_X1 _25758_ (.A(_16038_),
    .B(_01010_),
    .Z(_16039_));
 BUF_X2 _25759_ (.A(_03738_),
    .Z(_16040_));
 MUX2_X1 _25760_ (.A(_01221_),
    .B(_16039_),
    .S(_16040_),
    .Z(_01071_));
 XOR2_X1 _25761_ (.A(_17164_),
    .B(_16999_),
    .Z(_16041_));
 XOR2_X2 _25762_ (.A(_12385_),
    .B(_12807_),
    .Z(_16042_));
 XNOR2_X1 _25763_ (.A(_16042_),
    .B(_12651_),
    .ZN(_16043_));
 XNOR2_X1 _25764_ (.A(_16043_),
    .B(_13017_),
    .ZN(_16044_));
 XNOR2_X1 _25765_ (.A(_16044_),
    .B(_17164_),
    .ZN(_16045_));
 MUX2_X1 _25766_ (.A(_16041_),
    .B(_16045_),
    .S(_15155_),
    .Z(_00686_));
 NAND2_X1 _25767_ (.A1(_15524_),
    .A2(_15531_),
    .ZN(_16046_));
 AND2_X1 _25768_ (.A1(_15798_),
    .A2(_15799_),
    .ZN(_16047_));
 AND4_X1 _25769_ (.A1(_16046_),
    .A2(_16047_),
    .A3(_16004_),
    .A4(_15706_),
    .ZN(_16048_));
 OAI211_X1 _25770_ (.A(_15569_),
    .B(_15534_),
    .C1(_15475_),
    .C2(_15415_),
    .ZN(_16049_));
 AND4_X1 _25771_ (.A1(_15839_),
    .A2(_16049_),
    .A3(_15840_),
    .A4(_15841_),
    .ZN(_16050_));
 AND2_X1 _25772_ (.A1(_15569_),
    .A2(_15520_),
    .ZN(_16051_));
 AOI211_X1 _25773_ (.A(_16051_),
    .B(_15917_),
    .C1(_15570_),
    .C2(_15627_),
    .ZN(_16052_));
 AND2_X1 _25774_ (.A1(_15564_),
    .A2(_15498_),
    .ZN(_16053_));
 AND2_X1 _25775_ (.A1(_15498_),
    .A2(_15548_),
    .ZN(_16054_));
 OR4_X1 _25776_ (.A1(_15521_),
    .A2(_16053_),
    .A3(_15856_),
    .A4(_16054_),
    .ZN(_16055_));
 AND2_X1 _25777_ (.A1(_15444_),
    .A2(_15562_),
    .ZN(_16056_));
 AOI21_X1 _25778_ (.A(_15820_),
    .B1(_15732_),
    .B2(_15539_),
    .ZN(_16057_));
 NOR4_X1 _25779_ (.A1(_16055_),
    .A2(_16056_),
    .A3(_15924_),
    .A4(_16057_),
    .ZN(_16058_));
 AND4_X1 _25780_ (.A1(_16048_),
    .A2(_16050_),
    .A3(_16052_),
    .A4(_16058_),
    .ZN(_16059_));
 OAI21_X1 _25781_ (.A(_15512_),
    .B1(_15646_),
    .B2(_15516_),
    .ZN(_16060_));
 NAND3_X1 _25782_ (.A1(_15562_),
    .A2(_15429_),
    .A3(_15614_),
    .ZN(_16061_));
 OAI211_X1 _25783_ (.A(_16060_),
    .B(_16061_),
    .C1(_15763_),
    .C2(_15821_),
    .ZN(_16062_));
 AOI21_X1 _25784_ (.A(_15763_),
    .B1(_15631_),
    .B2(_15553_),
    .ZN(_16063_));
 AND4_X1 _25785_ (.A1(_15512_),
    .A2(_15460_),
    .A3(_15559_),
    .A4(_15534_),
    .ZN(_16064_));
 NOR3_X1 _25786_ (.A1(_16062_),
    .A2(_16063_),
    .A3(_16064_),
    .ZN(_16065_));
 NAND2_X1 _25787_ (.A1(_15588_),
    .A2(_15434_),
    .ZN(_16066_));
 NAND2_X1 _25788_ (.A1(_15886_),
    .A2(_16066_),
    .ZN(_16067_));
 AOI211_X1 _25789_ (.A(_16029_),
    .B(_16067_),
    .C1(_15602_),
    .C2(_15588_),
    .ZN(_16068_));
 AND2_X1 _25790_ (.A1(_15633_),
    .A2(_15507_),
    .ZN(_16069_));
 NAND2_X1 _25791_ (.A1(_15507_),
    .A2(_15520_),
    .ZN(_16070_));
 OAI21_X1 _25792_ (.A(_16070_),
    .B1(_15737_),
    .B2(_15555_),
    .ZN(_16071_));
 AND4_X1 _25793_ (.A1(_15436_),
    .A2(_15614_),
    .A3(_15534_),
    .A4(_15469_),
    .ZN(_16072_));
 AND4_X1 _25794_ (.A1(_15436_),
    .A2(_15614_),
    .A3(_15463_),
    .A4(_15469_),
    .ZN(_16073_));
 NOR4_X1 _25795_ (.A1(_16069_),
    .A2(_16071_),
    .A3(_16072_),
    .A4(_16073_),
    .ZN(_16074_));
 AOI21_X1 _25796_ (.A(_15881_),
    .B1(_15537_),
    .B2(_15632_),
    .ZN(_16075_));
 AOI211_X1 _25797_ (.A(_15743_),
    .B(_16075_),
    .C1(_15611_),
    .C2(_15797_),
    .ZN(_16076_));
 AND4_X1 _25798_ (.A1(_16065_),
    .A2(_16068_),
    .A3(_16074_),
    .A4(_16076_),
    .ZN(_16077_));
 OAI21_X1 _25799_ (.A(_15523_),
    .B1(_15527_),
    .B2(_15572_),
    .ZN(_16078_));
 OAI21_X1 _25800_ (.A(_15523_),
    .B1(_15849_),
    .B2(_15646_),
    .ZN(_16079_));
 AND2_X1 _25801_ (.A1(_16078_),
    .A2(_16079_),
    .ZN(_16080_));
 AND2_X1 _25802_ (.A1(_15412_),
    .A2(_15516_),
    .ZN(_16081_));
 NAND2_X1 _25803_ (.A1(_15412_),
    .A2(_15552_),
    .ZN(_16082_));
 NAND2_X1 _25804_ (.A1(_15412_),
    .A2(_15456_),
    .ZN(_16083_));
 OAI221_X1 _25805_ (.A(_16082_),
    .B1(_15544_),
    .B2(_15543_),
    .C1(_15436_),
    .C2(_16083_),
    .ZN(_16084_));
 AOI211_X1 _25806_ (.A(_16081_),
    .B(_16084_),
    .C1(_15413_),
    .C2(_15602_),
    .ZN(_16085_));
 AND2_X1 _25807_ (.A1(_15545_),
    .A2(_15578_),
    .ZN(_16086_));
 NOR4_X1 _25808_ (.A1(_15600_),
    .A2(_15653_),
    .A3(_16086_),
    .A4(_15862_),
    .ZN(_16087_));
 AND2_X1 _25809_ (.A1(_15430_),
    .A2(_15605_),
    .ZN(_16088_));
 OAI21_X1 _25810_ (.A(_15671_),
    .B1(_15683_),
    .B2(_15848_),
    .ZN(_16089_));
 AOI211_X1 _25811_ (.A(_16088_),
    .B(_16089_),
    .C1(_15654_),
    .C2(_15431_),
    .ZN(_16090_));
 AND4_X1 _25812_ (.A1(_16080_),
    .A2(_16085_),
    .A3(_16087_),
    .A4(_16090_),
    .ZN(_16091_));
 OAI21_X1 _25813_ (.A(_15618_),
    .B1(_15849_),
    .B2(_15646_),
    .ZN(_16092_));
 OAI21_X1 _25814_ (.A(_15453_),
    .B1(_15419_),
    .B2(_15434_),
    .ZN(_16093_));
 NAND4_X1 _25815_ (.A1(_15449_),
    .A2(_15534_),
    .A3(_15436_),
    .A4(_15451_),
    .ZN(_16094_));
 AND3_X1 _25816_ (.A1(_16092_),
    .A2(_16093_),
    .A3(_16094_),
    .ZN(_16095_));
 AOI21_X1 _25817_ (.A(_15786_),
    .B1(_15567_),
    .B2(_15851_),
    .ZN(_16096_));
 AOI211_X1 _25818_ (.A(_15594_),
    .B(_15786_),
    .C1(_15599_),
    .C2(_15559_),
    .ZN(_16097_));
 AOI211_X1 _25819_ (.A(_16096_),
    .B(_16097_),
    .C1(_15572_),
    .C2(_15637_),
    .ZN(_16098_));
 AOI21_X1 _25820_ (.A(_15674_),
    .B1(_15732_),
    .B2(_15918_),
    .ZN(_16099_));
 AND2_X1 _25821_ (.A1(_15690_),
    .A2(_15470_),
    .ZN(_16100_));
 AND2_X1 _25822_ (.A1(_15652_),
    .A2(_15470_),
    .ZN(_16101_));
 NOR4_X1 _25823_ (.A1(_16099_),
    .A2(_16100_),
    .A3(_16101_),
    .A4(_15679_),
    .ZN(_16102_));
 NOR2_X1 _25824_ (.A1(_15783_),
    .A2(_15692_),
    .ZN(_16103_));
 NAND2_X1 _25825_ (.A1(_15565_),
    .A2(_15484_),
    .ZN(_16104_));
 AND2_X1 _25826_ (.A1(_15484_),
    .A2(_15551_),
    .ZN(_16105_));
 INV_X1 _25827_ (.A(_16105_),
    .ZN(_16106_));
 AND4_X1 _25828_ (.A1(_15621_),
    .A2(_16103_),
    .A3(_16104_),
    .A4(_16106_),
    .ZN(_16107_));
 AND4_X1 _25829_ (.A1(_16095_),
    .A2(_16098_),
    .A3(_16102_),
    .A4(_16107_),
    .ZN(_16108_));
 NAND4_X1 _25830_ (.A1(_16059_),
    .A2(_16077_),
    .A3(_16091_),
    .A4(_16108_),
    .ZN(_16109_));
 NOR2_X1 _25831_ (.A1(_16109_),
    .A2(_15575_),
    .ZN(_16110_));
 INV_X1 _25832_ (.A(_01011_),
    .ZN(_16111_));
 XNOR2_X1 _25833_ (.A(_16110_),
    .B(_16111_),
    .ZN(_16112_));
 MUX2_X1 _25834_ (.A(_01222_),
    .B(_16112_),
    .S(_16040_),
    .Z(_01072_));
 OR4_X1 _25835_ (.A1(_15448_),
    .A2(_15826_),
    .A3(_15858_),
    .A4(_15468_),
    .ZN(_16113_));
 OAI211_X1 _25836_ (.A(_15499_),
    .B(_15473_),
    .C1(_15459_),
    .C2(_15486_),
    .ZN(_16114_));
 OAI21_X1 _25837_ (.A(_16114_),
    .B1(_15789_),
    .B2(_15556_),
    .ZN(_16115_));
 NOR4_X1 _25838_ (.A1(_16113_),
    .A2(_15723_),
    .A3(_16054_),
    .A4(_16115_),
    .ZN(_16116_));
 OAI211_X1 _25839_ (.A(_16015_),
    .B(_15671_),
    .C1(_15683_),
    .C2(_15848_),
    .ZN(_16117_));
 INV_X1 _25840_ (.A(_15814_),
    .ZN(_16118_));
 OAI21_X1 _25841_ (.A(_15413_),
    .B1(_15592_),
    .B2(_15440_),
    .ZN(_16119_));
 NAND4_X1 _25842_ (.A1(_16118_),
    .A2(_16083_),
    .A3(_16082_),
    .A4(_16119_),
    .ZN(_16120_));
 OAI21_X1 _25843_ (.A(_15947_),
    .B1(_15918_),
    .B2(_15848_),
    .ZN(_16121_));
 NOR4_X1 _25844_ (.A1(_16117_),
    .A2(_16120_),
    .A3(_15549_),
    .A4(_16121_),
    .ZN(_16122_));
 INV_X1 _25845_ (.A(_16000_),
    .ZN(_16123_));
 AOI211_X1 _25846_ (.A(_15712_),
    .B(_15835_),
    .C1(_15532_),
    .C2(_15854_),
    .ZN(_16124_));
 OAI21_X1 _25847_ (.A(_15570_),
    .B1(_15797_),
    .B2(_15533_),
    .ZN(_16125_));
 OAI21_X1 _25848_ (.A(_15570_),
    .B1(_15493_),
    .B2(_15552_),
    .ZN(_16126_));
 AND4_X1 _25849_ (.A1(_16123_),
    .A2(_16124_),
    .A3(_16125_),
    .A4(_16126_),
    .ZN(_16127_));
 AOI21_X1 _25850_ (.A(_15546_),
    .B1(_15880_),
    .B2(_15927_),
    .ZN(_16128_));
 OAI211_X1 _25851_ (.A(_15932_),
    .B(_16009_),
    .C1(_15650_),
    .C2(_15546_),
    .ZN(_16129_));
 AOI21_X1 _25852_ (.A(_15550_),
    .B1(_15732_),
    .B2(_15918_),
    .ZN(_16130_));
 AOI21_X1 _25853_ (.A(_15550_),
    .B1(_15789_),
    .B2(_15790_),
    .ZN(_16131_));
 NOR4_X1 _25854_ (.A1(_16128_),
    .A2(_16129_),
    .A3(_16130_),
    .A4(_16131_),
    .ZN(_16132_));
 NAND4_X1 _25855_ (.A1(_16116_),
    .A2(_16122_),
    .A3(_16127_),
    .A4(_16132_),
    .ZN(_16133_));
 AOI22_X1 _25856_ (.A1(_15777_),
    .A2(_15460_),
    .B1(_15434_),
    .B2(_15471_),
    .ZN(_16134_));
 AND2_X1 _25857_ (.A1(_15618_),
    .A2(_15520_),
    .ZN(_16135_));
 AND2_X1 _25858_ (.A1(_15565_),
    .A2(_15618_),
    .ZN(_16136_));
 AOI211_X1 _25859_ (.A(_16135_),
    .B(_16136_),
    .C1(_15554_),
    .C2(_15618_),
    .ZN(_16137_));
 NOR3_X1 _25860_ (.A1(_15773_),
    .A2(_16101_),
    .A3(_15680_),
    .ZN(_16138_));
 OAI211_X1 _25861_ (.A(_15618_),
    .B(_15486_),
    .C1(_15598_),
    .C2(_15535_),
    .ZN(_16139_));
 AND4_X1 _25862_ (.A1(_16134_),
    .A2(_16137_),
    .A3(_16138_),
    .A4(_16139_),
    .ZN(_16140_));
 NAND2_X1 _25863_ (.A1(_15604_),
    .A2(_15652_),
    .ZN(_16141_));
 AOI21_X1 _25864_ (.A(_15882_),
    .B1(_15611_),
    .B2(_16023_),
    .ZN(_16142_));
 OAI21_X1 _25865_ (.A(_15604_),
    .B1(_15633_),
    .B2(_15572_),
    .ZN(_16143_));
 OAI21_X1 _25866_ (.A(_15611_),
    .B1(_15524_),
    .B2(_15548_),
    .ZN(_16144_));
 AND4_X1 _25867_ (.A1(_16141_),
    .A2(_16142_),
    .A3(_16143_),
    .A4(_16144_),
    .ZN(_16145_));
 AND3_X1 _25868_ (.A1(_15694_),
    .A2(_15487_),
    .A3(_15488_),
    .ZN(_16146_));
 AND2_X1 _25869_ (.A1(_15572_),
    .A2(_15485_),
    .ZN(_16147_));
 AND2_X1 _25870_ (.A1(_15493_),
    .A2(_15484_),
    .ZN(_16148_));
 NOR4_X1 _25871_ (.A1(_16147_),
    .A2(_15788_),
    .A3(_16148_),
    .A4(_16105_),
    .ZN(_16149_));
 AND2_X1 _25872_ (.A1(_15447_),
    .A2(_15637_),
    .ZN(_16150_));
 AND2_X1 _25873_ (.A1(_15637_),
    .A2(_15865_),
    .ZN(_16151_));
 NOR4_X1 _25874_ (.A1(_15702_),
    .A2(_15951_),
    .A3(_16150_),
    .A4(_16151_),
    .ZN(_16152_));
 AND3_X1 _25875_ (.A1(_16146_),
    .A2(_16149_),
    .A3(_16152_),
    .ZN(_16153_));
 NAND2_X1 _25876_ (.A1(_15627_),
    .A2(_15513_),
    .ZN(_16154_));
 AND2_X1 _25877_ (.A1(_16154_),
    .A2(_16061_),
    .ZN(_16155_));
 OAI221_X1 _25878_ (.A(_15588_),
    .B1(_15437_),
    .B2(_10946_),
    .C1(_15473_),
    .C2(_15464_),
    .ZN(_16156_));
 OAI21_X1 _25879_ (.A(_15513_),
    .B1(_15595_),
    .B2(_15552_),
    .ZN(_16157_));
 AND4_X1 _25880_ (.A1(_16155_),
    .A2(_16066_),
    .A3(_16156_),
    .A4(_16157_),
    .ZN(_16158_));
 NAND4_X1 _25881_ (.A1(_16140_),
    .A2(_16145_),
    .A3(_16153_),
    .A4(_16158_),
    .ZN(_16159_));
 NOR2_X1 _25882_ (.A1(_16133_),
    .A2(_16159_),
    .ZN(_16160_));
 XOR2_X1 _25883_ (.A(_16160_),
    .B(_01012_),
    .Z(_16161_));
 MUX2_X1 _25884_ (.A(_01223_),
    .B(_16161_),
    .S(_16040_),
    .Z(_01073_));
 INV_X1 _25885_ (.A(_17074_),
    .ZN(_16162_));
 NOR2_X2 _25886_ (.A1(_16162_),
    .A2(_17075_),
    .ZN(_16163_));
 BUF_X2 _25887_ (.A(_16163_),
    .Z(_16164_));
 INV_X1 _25888_ (.A(_16164_),
    .ZN(_16165_));
 NOR2_X2 _25889_ (.A1(_11012_),
    .A2(_17076_),
    .ZN(_16166_));
 CLKBUF_X2 _25890_ (.A(_16166_),
    .Z(_16167_));
 NAND2_X1 _25891_ (.A1(_16165_),
    .A2(_16167_),
    .ZN(_16168_));
 INV_X1 _25892_ (.A(_17075_),
    .ZN(_16169_));
 NOR2_X2 _25893_ (.A1(_16169_),
    .A2(_17074_),
    .ZN(_16170_));
 CLKBUF_X2 _25894_ (.A(_16170_),
    .Z(_16171_));
 NOR2_X1 _25895_ (.A1(_16168_),
    .A2(_16171_),
    .ZN(_16172_));
 INV_X1 _25896_ (.A(_17080_),
    .ZN(_16173_));
 AND2_X1 _25897_ (.A1(_16173_),
    .A2(_17079_),
    .ZN(_16174_));
 CLKBUF_X2 _25898_ (.A(_16174_),
    .Z(_16175_));
 NOR2_X2 _25899_ (.A1(_17081_),
    .A2(_17082_),
    .ZN(_16176_));
 AND2_X1 _25900_ (.A1(_16175_),
    .A2(_16176_),
    .ZN(_16177_));
 BUF_X2 _25901_ (.A(_16177_),
    .Z(_16178_));
 NAND2_X1 _25902_ (.A1(_16172_),
    .A2(_16178_),
    .ZN(_16179_));
 BUF_X2 _25903_ (.A(_16178_),
    .Z(_16180_));
 NOR2_X1 _25904_ (.A1(_17076_),
    .A2(_17077_),
    .ZN(_16181_));
 CLKBUF_X2 _25905_ (.A(_16181_),
    .Z(_16182_));
 AND2_X2 _25906_ (.A1(_16182_),
    .A2(_17075_),
    .ZN(_16183_));
 NAND2_X1 _25907_ (.A1(_16180_),
    .A2(_16183_),
    .ZN(_16184_));
 INV_X1 _25908_ (.A(_16178_),
    .ZN(_16185_));
 NOR2_X2 _25909_ (.A1(_17074_),
    .A2(_17075_),
    .ZN(_16186_));
 INV_X2 _25910_ (.A(_16186_),
    .ZN(_16187_));
 INV_X1 _25911_ (.A(_17076_),
    .ZN(_16188_));
 NOR2_X2 _25912_ (.A1(_16188_),
    .A2(_17077_),
    .ZN(_16189_));
 CLKBUF_X2 _25913_ (.A(_16189_),
    .Z(_16190_));
 NAND2_X1 _25914_ (.A1(_16187_),
    .A2(_16190_),
    .ZN(_16191_));
 AND2_X1 _25915_ (.A1(_17074_),
    .A2(_17075_),
    .ZN(_16192_));
 BUF_X2 _25916_ (.A(_16192_),
    .Z(_16193_));
 NOR2_X1 _25917_ (.A1(_16191_),
    .A2(_16193_),
    .ZN(_16194_));
 INV_X1 _25918_ (.A(_16194_),
    .ZN(_16195_));
 OAI211_X1 _25919_ (.A(_16179_),
    .B(_16184_),
    .C1(_16185_),
    .C2(_16195_),
    .ZN(_16196_));
 AND2_X2 _25920_ (.A1(_16189_),
    .A2(_17075_),
    .ZN(_16197_));
 NOR2_X1 _25921_ (.A1(_17079_),
    .A2(_17080_),
    .ZN(_16198_));
 AND2_X1 _25922_ (.A1(_16198_),
    .A2(_16176_),
    .ZN(_16199_));
 AND2_X1 _25923_ (.A1(_16197_),
    .A2(_16199_),
    .ZN(_16200_));
 INV_X1 _25924_ (.A(_16200_),
    .ZN(_16201_));
 NAND3_X1 _25925_ (.A1(_16199_),
    .A2(_16190_),
    .A3(_16164_),
    .ZN(_16202_));
 INV_X1 _25926_ (.A(_16183_),
    .ZN(_16203_));
 INV_X1 _25927_ (.A(_16199_),
    .ZN(_16204_));
 OAI211_X1 _25928_ (.A(_16201_),
    .B(_16202_),
    .C1(_16203_),
    .C2(_16204_),
    .ZN(_16205_));
 AND2_X1 _25929_ (.A1(_16166_),
    .A2(_17075_),
    .ZN(_16206_));
 BUF_X2 _25930_ (.A(_16206_),
    .Z(_16207_));
 NAND2_X1 _25931_ (.A1(_16207_),
    .A2(_16199_),
    .ZN(_16208_));
 NAND3_X1 _25932_ (.A1(_16199_),
    .A2(_16164_),
    .A3(_16167_),
    .ZN(_16209_));
 AND2_X1 _25933_ (.A1(_17076_),
    .A2(_17077_),
    .ZN(_16210_));
 AND2_X1 _25934_ (.A1(_16170_),
    .A2(_16210_),
    .ZN(_16211_));
 AND2_X1 _25935_ (.A1(_16163_),
    .A2(_16210_),
    .ZN(_16212_));
 NOR2_X1 _25936_ (.A1(_16211_),
    .A2(_16212_),
    .ZN(_16213_));
 OAI211_X1 _25937_ (.A(_16208_),
    .B(_16209_),
    .C1(_16213_),
    .C2(_16204_),
    .ZN(_16214_));
 NOR3_X1 _25938_ (.A1(_16196_),
    .A2(_16205_),
    .A3(_16214_),
    .ZN(_16215_));
 INV_X1 _25939_ (.A(_16193_),
    .ZN(_16216_));
 NOR2_X1 _25940_ (.A1(_16173_),
    .A2(_17079_),
    .ZN(_16217_));
 AND2_X2 _25941_ (.A1(_16217_),
    .A2(_16176_),
    .ZN(_16218_));
 BUF_X2 _25942_ (.A(_16218_),
    .Z(_16219_));
 INV_X1 _25943_ (.A(_16191_),
    .ZN(_16220_));
 BUF_X2 _25944_ (.A(_16182_),
    .Z(_16221_));
 OAI211_X1 _25945_ (.A(_16216_),
    .B(_16219_),
    .C1(_16220_),
    .C2(_16221_),
    .ZN(_16222_));
 CLKBUF_X2 _25946_ (.A(_16210_),
    .Z(_16223_));
 AND2_X1 _25947_ (.A1(_16223_),
    .A2(_16186_),
    .ZN(_16224_));
 CLKBUF_X2 _25948_ (.A(_16217_),
    .Z(_16225_));
 AND3_X1 _25949_ (.A1(_16224_),
    .A2(_16225_),
    .A3(_16176_),
    .ZN(_16226_));
 AND2_X1 _25950_ (.A1(_16223_),
    .A2(_17075_),
    .ZN(_16227_));
 CLKBUF_X2 _25951_ (.A(_16227_),
    .Z(_16228_));
 AND2_X1 _25952_ (.A1(_16218_),
    .A2(_16228_),
    .ZN(_16229_));
 BUF_X2 _25953_ (.A(_16167_),
    .Z(_16230_));
 NAND2_X1 _25954_ (.A1(_16187_),
    .A2(_16230_),
    .ZN(_16231_));
 INV_X1 _25955_ (.A(_16231_),
    .ZN(_16232_));
 AOI211_X1 _25956_ (.A(_16226_),
    .B(_16229_),
    .C1(_16219_),
    .C2(_16232_),
    .ZN(_16233_));
 INV_X1 _25957_ (.A(_16223_),
    .ZN(_16234_));
 AND2_X1 _25958_ (.A1(_17079_),
    .A2(_17080_),
    .ZN(_16235_));
 CLKBUF_X2 _25959_ (.A(_16235_),
    .Z(_16236_));
 AND2_X2 _25960_ (.A1(_16236_),
    .A2(_16176_),
    .ZN(_16237_));
 INV_X1 _25961_ (.A(_16237_),
    .ZN(_16238_));
 BUF_X2 _25962_ (.A(_16162_),
    .Z(_16239_));
 AOI211_X1 _25963_ (.A(_16234_),
    .B(_16238_),
    .C1(_16239_),
    .C2(_10993_),
    .ZN(_16240_));
 AND3_X1 _25964_ (.A1(_16237_),
    .A2(_16190_),
    .A3(_16171_),
    .ZN(_16241_));
 NAND2_X1 _25965_ (.A1(_16187_),
    .A2(_16182_),
    .ZN(_16242_));
 NOR2_X1 _25966_ (.A1(_16238_),
    .A2(_16242_),
    .ZN(_16243_));
 AND2_X2 _25967_ (.A1(_16166_),
    .A2(_16186_),
    .ZN(_16244_));
 AND2_X1 _25968_ (.A1(_16244_),
    .A2(_16237_),
    .ZN(_16245_));
 NOR4_X1 _25969_ (.A1(_16240_),
    .A2(_16241_),
    .A3(_16243_),
    .A4(_16245_),
    .ZN(_16246_));
 AND4_X1 _25970_ (.A1(_16215_),
    .A2(_16222_),
    .A3(_16233_),
    .A4(_16246_),
    .ZN(_16247_));
 INV_X1 _25971_ (.A(_17081_),
    .ZN(_16248_));
 AND2_X1 _25972_ (.A1(_16248_),
    .A2(_17082_),
    .ZN(_16249_));
 AND2_X1 _25973_ (.A1(_16249_),
    .A2(_16198_),
    .ZN(_16250_));
 INV_X1 _25974_ (.A(_16250_),
    .ZN(_16251_));
 OR2_X1 _25975_ (.A1(_16213_),
    .A2(_16251_),
    .ZN(_16252_));
 AND2_X1 _25976_ (.A1(_16210_),
    .A2(_16192_),
    .ZN(_16253_));
 AND2_X1 _25977_ (.A1(_16250_),
    .A2(_16253_),
    .ZN(_16254_));
 INV_X1 _25978_ (.A(_16254_),
    .ZN(_16255_));
 NAND2_X1 _25979_ (.A1(_16252_),
    .A2(_16255_),
    .ZN(_16256_));
 AND2_X1 _25980_ (.A1(_16166_),
    .A2(_17074_),
    .ZN(_16257_));
 BUF_X2 _25981_ (.A(_16250_),
    .Z(_16258_));
 AOI21_X1 _25982_ (.A(_16256_),
    .B1(_16257_),
    .B2(_16258_),
    .ZN(_16259_));
 INV_X1 _25983_ (.A(_16190_),
    .ZN(_16260_));
 NOR2_X1 _25984_ (.A1(_16260_),
    .A2(_16170_),
    .ZN(_16261_));
 NAND2_X1 _25985_ (.A1(_16261_),
    .A2(_16250_),
    .ZN(_16262_));
 AND2_X1 _25986_ (.A1(_16175_),
    .A2(_16249_),
    .ZN(_16263_));
 CLKBUF_X2 _25987_ (.A(_16263_),
    .Z(_16264_));
 NOR3_X1 _25988_ (.A1(_16193_),
    .A2(_17076_),
    .A3(_17077_),
    .ZN(_16265_));
 AND3_X1 _25989_ (.A1(_16264_),
    .A2(_16187_),
    .A3(_16265_),
    .ZN(_16266_));
 AOI21_X1 _25990_ (.A(_16266_),
    .B1(_16228_),
    .B2(_16264_),
    .ZN(_16267_));
 BUF_X2 _25991_ (.A(_16249_),
    .Z(_16268_));
 BUF_X2 _25992_ (.A(_16268_),
    .Z(_16269_));
 BUF_X2 _25993_ (.A(_16198_),
    .Z(_16270_));
 NAND4_X1 _25994_ (.A1(_16269_),
    .A2(_16239_),
    .A3(_16221_),
    .A4(_16270_),
    .ZN(_16271_));
 NAND4_X1 _25995_ (.A1(_16259_),
    .A2(_16262_),
    .A3(_16267_),
    .A4(_16271_),
    .ZN(_16272_));
 AND2_X1 _25996_ (.A1(_16189_),
    .A2(_16186_),
    .ZN(_16273_));
 AND3_X1 _25997_ (.A1(_16273_),
    .A2(_16217_),
    .A3(_16249_),
    .ZN(_16274_));
 BUF_X2 _25998_ (.A(_16253_),
    .Z(_16275_));
 BUF_X2 _25999_ (.A(_16169_),
    .Z(_16276_));
 AND2_X1 _26000_ (.A1(_16223_),
    .A2(_16276_),
    .ZN(_16277_));
 CLKBUF_X2 _26001_ (.A(_16277_),
    .Z(_16278_));
 OAI211_X1 _26002_ (.A(_16225_),
    .B(_16269_),
    .C1(_16275_),
    .C2(_16278_),
    .ZN(_16279_));
 AND2_X1 _26003_ (.A1(_16249_),
    .A2(_16217_),
    .ZN(_16280_));
 BUF_X2 _26004_ (.A(_16280_),
    .Z(_16281_));
 INV_X1 _26005_ (.A(_16281_),
    .ZN(_16282_));
 AND2_X2 _26006_ (.A1(_16163_),
    .A2(_16166_),
    .ZN(_16283_));
 INV_X1 _26007_ (.A(_16283_),
    .ZN(_16284_));
 OAI21_X1 _26008_ (.A(_16279_),
    .B1(_16282_),
    .B2(_16284_),
    .ZN(_16285_));
 AND2_X1 _26009_ (.A1(_16249_),
    .A2(_16235_),
    .ZN(_16286_));
 AND2_X1 _26010_ (.A1(_16261_),
    .A2(_16286_),
    .ZN(_16287_));
 AND2_X1 _26011_ (.A1(_16286_),
    .A2(_16224_),
    .ZN(_16288_));
 INV_X1 _26012_ (.A(_16182_),
    .ZN(_16289_));
 NOR2_X2 _26013_ (.A1(_16289_),
    .A2(_16163_),
    .ZN(_16290_));
 AND2_X1 _26014_ (.A1(_16286_),
    .A2(_16290_),
    .ZN(_16291_));
 OR3_X1 _26015_ (.A1(_16287_),
    .A2(_16288_),
    .A3(_16291_),
    .ZN(_16292_));
 NOR4_X1 _26016_ (.A1(_16272_),
    .A2(_16274_),
    .A3(_16285_),
    .A4(_16292_),
    .ZN(_16293_));
 AND2_X1 _26017_ (.A1(_17081_),
    .A2(_17082_),
    .ZN(_16294_));
 AND2_X2 _26018_ (.A1(_16217_),
    .A2(_16294_),
    .ZN(_16295_));
 CLKBUF_X2 _26019_ (.A(_16295_),
    .Z(_16296_));
 AND2_X1 _26020_ (.A1(_16192_),
    .A2(_16181_),
    .ZN(_16297_));
 INV_X1 _26021_ (.A(_16297_),
    .ZN(_16298_));
 AND2_X1 _26022_ (.A1(_16182_),
    .A2(_16186_),
    .ZN(_16299_));
 INV_X1 _26023_ (.A(_16299_),
    .ZN(_16300_));
 NAND2_X1 _26024_ (.A1(_16298_),
    .A2(_16300_),
    .ZN(_16301_));
 AND2_X2 _26025_ (.A1(_16189_),
    .A2(_16276_),
    .ZN(_16302_));
 OAI21_X1 _26026_ (.A(_16296_),
    .B1(_16301_),
    .B2(_16302_),
    .ZN(_16303_));
 AND2_X1 _26027_ (.A1(_16174_),
    .A2(_16294_),
    .ZN(_16304_));
 CLKBUF_X2 _26028_ (.A(_16304_),
    .Z(_16305_));
 AND2_X2 _26029_ (.A1(_16190_),
    .A2(_16164_),
    .ZN(_16306_));
 AND2_X1 _26030_ (.A1(_16170_),
    .A2(_16182_),
    .ZN(_16307_));
 CLKBUF_X2 _26031_ (.A(_16307_),
    .Z(_16308_));
 OAI21_X1 _26032_ (.A(_16305_),
    .B1(_16306_),
    .B2(_16308_),
    .ZN(_16309_));
 AND2_X1 _26033_ (.A1(_16166_),
    .A2(_16169_),
    .ZN(_16310_));
 AND2_X1 _26034_ (.A1(_16305_),
    .A2(_16310_),
    .ZN(_16311_));
 AND2_X1 _26035_ (.A1(_16166_),
    .A2(_16193_),
    .ZN(_16312_));
 AND2_X1 _26036_ (.A1(_16304_),
    .A2(_16312_),
    .ZN(_16313_));
 AND2_X1 _26037_ (.A1(_16170_),
    .A2(_16166_),
    .ZN(_16314_));
 BUF_X2 _26038_ (.A(_16314_),
    .Z(_16315_));
 AOI211_X1 _26039_ (.A(_16311_),
    .B(_16313_),
    .C1(_16305_),
    .C2(_16315_),
    .ZN(_16316_));
 BUF_X2 _26040_ (.A(_16211_),
    .Z(_16317_));
 CLKBUF_X2 _26041_ (.A(_16212_),
    .Z(_16318_));
 OAI21_X1 _26042_ (.A(_16305_),
    .B1(_16317_),
    .B2(_16318_),
    .ZN(_16319_));
 AND2_X1 _26043_ (.A1(_16294_),
    .A2(_16198_),
    .ZN(_16320_));
 NAND2_X1 _26044_ (.A1(_16212_),
    .A2(_16320_),
    .ZN(_16321_));
 CLKBUF_X2 _26045_ (.A(_16320_),
    .Z(_16322_));
 NAND2_X1 _26046_ (.A1(_16224_),
    .A2(_16322_),
    .ZN(_16323_));
 NAND2_X1 _26047_ (.A1(_16321_),
    .A2(_16323_),
    .ZN(_16324_));
 AND2_X1 _26048_ (.A1(_16257_),
    .A2(_16320_),
    .ZN(_16325_));
 AND2_X1 _26049_ (.A1(_16307_),
    .A2(_16320_),
    .ZN(_16326_));
 BUF_X2 _26050_ (.A(_16294_),
    .Z(_16327_));
 AND4_X1 _26051_ (.A1(_16327_),
    .A2(_16170_),
    .A3(_16223_),
    .A4(_16198_),
    .ZN(_16328_));
 NOR4_X1 _26052_ (.A1(_16324_),
    .A2(_16325_),
    .A3(_16326_),
    .A4(_16328_),
    .ZN(_16329_));
 AND4_X1 _26053_ (.A1(_16309_),
    .A2(_16316_),
    .A3(_16319_),
    .A4(_16329_),
    .ZN(_16330_));
 AND2_X1 _26054_ (.A1(_16223_),
    .A2(_10986_),
    .ZN(_16331_));
 AND2_X1 _26055_ (.A1(_16295_),
    .A2(_16331_),
    .ZN(_16332_));
 NAND2_X1 _26056_ (.A1(_16312_),
    .A2(_16295_),
    .ZN(_16333_));
 INV_X1 _26057_ (.A(_16315_),
    .ZN(_16334_));
 INV_X1 _26058_ (.A(_16295_),
    .ZN(_16335_));
 OAI21_X1 _26059_ (.A(_16333_),
    .B1(_16334_),
    .B2(_16335_),
    .ZN(_16336_));
 AOI211_X1 _26060_ (.A(_16332_),
    .B(_16336_),
    .C1(_16244_),
    .C2(_16296_),
    .ZN(_16337_));
 AND2_X1 _26061_ (.A1(_16294_),
    .A2(_16235_),
    .ZN(_16338_));
 CLKBUF_X2 _26062_ (.A(_16338_),
    .Z(_16339_));
 AND2_X1 _26063_ (.A1(_16317_),
    .A2(_16339_),
    .ZN(_16340_));
 AND2_X1 _26064_ (.A1(_16273_),
    .A2(_16338_),
    .ZN(_16341_));
 INV_X1 _26065_ (.A(_16341_),
    .ZN(_16342_));
 AND2_X1 _26066_ (.A1(_16163_),
    .A2(_16182_),
    .ZN(_16343_));
 BUF_X2 _26067_ (.A(_16343_),
    .Z(_16344_));
 NAND2_X1 _26068_ (.A1(_16344_),
    .A2(_16339_),
    .ZN(_16345_));
 INV_X1 _26069_ (.A(_16339_),
    .ZN(_16346_));
 OAI211_X1 _26070_ (.A(_16342_),
    .B(_16345_),
    .C1(_16203_),
    .C2(_16346_),
    .ZN(_16347_));
 CLKBUF_X2 _26071_ (.A(_16339_),
    .Z(_16348_));
 AOI211_X1 _26072_ (.A(_16340_),
    .B(_16347_),
    .C1(_16230_),
    .C2(_16348_),
    .ZN(_16349_));
 AND4_X1 _26073_ (.A1(_16303_),
    .A2(_16330_),
    .A3(_16337_),
    .A4(_16349_),
    .ZN(_16350_));
 NOR2_X1 _26074_ (.A1(_16248_),
    .A2(_17082_),
    .ZN(_16351_));
 AND2_X1 _26075_ (.A1(_16217_),
    .A2(_16351_),
    .ZN(_16352_));
 AND2_X1 _26076_ (.A1(_16352_),
    .A2(_16211_),
    .ZN(_16353_));
 AND2_X2 _26077_ (.A1(_16189_),
    .A2(_16170_),
    .ZN(_16354_));
 AND2_X1 _26078_ (.A1(_16352_),
    .A2(_16354_),
    .ZN(_16355_));
 INV_X1 _26079_ (.A(_16355_),
    .ZN(_16356_));
 AND2_X2 _26080_ (.A1(_16189_),
    .A2(_16193_),
    .ZN(_16357_));
 AND2_X1 _26081_ (.A1(_16352_),
    .A2(_16357_),
    .ZN(_16358_));
 INV_X1 _26082_ (.A(_16358_),
    .ZN(_16359_));
 BUF_X2 _26083_ (.A(_16352_),
    .Z(_16360_));
 NAND2_X1 _26084_ (.A1(_16360_),
    .A2(_16302_),
    .ZN(_16361_));
 NAND3_X1 _26085_ (.A1(_16356_),
    .A2(_16359_),
    .A3(_16361_),
    .ZN(_16362_));
 NAND2_X1 _26086_ (.A1(_16360_),
    .A2(_16344_),
    .ZN(_16363_));
 NAND2_X1 _26087_ (.A1(_16360_),
    .A2(_16297_),
    .ZN(_16364_));
 NAND2_X1 _26088_ (.A1(_16363_),
    .A2(_16364_),
    .ZN(_16365_));
 NAND2_X1 _26089_ (.A1(_16352_),
    .A2(_16312_),
    .ZN(_16366_));
 CLKBUF_X2 _26090_ (.A(_16351_),
    .Z(_16367_));
 NAND4_X1 _26091_ (.A1(_16167_),
    .A2(_16225_),
    .A3(_16367_),
    .A4(_16276_),
    .ZN(_16368_));
 NAND2_X1 _26092_ (.A1(_16366_),
    .A2(_16368_),
    .ZN(_16369_));
 OR4_X1 _26093_ (.A1(_16353_),
    .A2(_16362_),
    .A3(_16365_),
    .A4(_16369_),
    .ZN(_16370_));
 AND2_X1 _26094_ (.A1(_16367_),
    .A2(_16198_),
    .ZN(_16371_));
 OAI21_X1 _26095_ (.A(_16371_),
    .B1(_16317_),
    .B2(_16277_),
    .ZN(_16372_));
 NAND4_X1 _26096_ (.A1(_16167_),
    .A2(_16367_),
    .A3(_10986_),
    .A4(_16270_),
    .ZN(_16373_));
 AND2_X1 _26097_ (.A1(_16372_),
    .A2(_16373_),
    .ZN(_16374_));
 BUF_X2 _26098_ (.A(_16371_),
    .Z(_16375_));
 NAND2_X1 _26099_ (.A1(_16273_),
    .A2(_16375_),
    .ZN(_16376_));
 AND2_X2 _26100_ (.A1(_16182_),
    .A2(_16276_),
    .ZN(_16377_));
 INV_X1 _26101_ (.A(_16377_),
    .ZN(_16378_));
 INV_X1 _26102_ (.A(_16371_),
    .ZN(_16379_));
 OAI211_X1 _26103_ (.A(_16374_),
    .B(_16376_),
    .C1(_16378_),
    .C2(_16379_),
    .ZN(_16380_));
 AND2_X2 _26104_ (.A1(_16175_),
    .A2(_16351_),
    .ZN(_16381_));
 AND2_X1 _26105_ (.A1(_16381_),
    .A2(_16297_),
    .ZN(_16382_));
 AND2_X1 _26106_ (.A1(_16381_),
    .A2(_16377_),
    .ZN(_16383_));
 NOR2_X1 _26107_ (.A1(_16382_),
    .A2(_16383_),
    .ZN(_16384_));
 BUF_X2 _26108_ (.A(_16381_),
    .Z(_16385_));
 NAND2_X1 _26109_ (.A1(_16385_),
    .A2(_16197_),
    .ZN(_16386_));
 OAI21_X1 _26110_ (.A(_16385_),
    .B1(_16257_),
    .B2(_16275_),
    .ZN(_16387_));
 NAND3_X1 _26111_ (.A1(_16384_),
    .A2(_16386_),
    .A3(_16387_),
    .ZN(_16388_));
 NOR2_X1 _26112_ (.A1(_16211_),
    .A2(_16312_),
    .ZN(_16389_));
 AND2_X1 _26113_ (.A1(_16351_),
    .A2(_16236_),
    .ZN(_16390_));
 INV_X1 _26114_ (.A(_16390_),
    .ZN(_16391_));
 NOR2_X1 _26115_ (.A1(_16389_),
    .A2(_16391_),
    .ZN(_16392_));
 AND2_X1 _26116_ (.A1(_16212_),
    .A2(_16390_),
    .ZN(_16393_));
 NOR2_X1 _26117_ (.A1(_16392_),
    .A2(_16393_),
    .ZN(_16394_));
 NAND3_X1 _26118_ (.A1(_16377_),
    .A2(_16236_),
    .A3(_16367_),
    .ZN(_16395_));
 CLKBUF_X2 _26119_ (.A(_16390_),
    .Z(_16396_));
 BUF_X2 _26120_ (.A(_16297_),
    .Z(_16397_));
 NAND2_X1 _26121_ (.A1(_16396_),
    .A2(_16397_),
    .ZN(_16398_));
 AND2_X1 _26122_ (.A1(_16190_),
    .A2(_10986_),
    .ZN(_16399_));
 NAND2_X1 _26123_ (.A1(_16399_),
    .A2(_16396_),
    .ZN(_16400_));
 NAND4_X1 _26124_ (.A1(_16394_),
    .A2(_16395_),
    .A3(_16398_),
    .A4(_16400_),
    .ZN(_16401_));
 NOR4_X1 _26125_ (.A1(_16370_),
    .A2(_16380_),
    .A3(_16388_),
    .A4(_16401_),
    .ZN(_16402_));
 AND4_X1 _26126_ (.A1(_16247_),
    .A2(_16293_),
    .A3(_16350_),
    .A4(_16402_),
    .ZN(_16403_));
 OAI21_X1 _26127_ (.A(_11012_),
    .B1(_16187_),
    .B2(_17076_),
    .ZN(_16404_));
 AND3_X1 _26128_ (.A1(_16270_),
    .A2(_16176_),
    .A3(_11012_),
    .ZN(_16405_));
 AND2_X1 _26129_ (.A1(_16404_),
    .A2(_16405_),
    .ZN(_16406_));
 INV_X1 _26130_ (.A(_16406_),
    .ZN(_16407_));
 NAND2_X1 _26131_ (.A1(_16403_),
    .A2(_16407_),
    .ZN(_16408_));
 XNOR2_X1 _26132_ (.A(_01014_),
    .B(_01013_),
    .ZN(_16409_));
 XNOR2_X1 _26133_ (.A(_16408_),
    .B(_16409_),
    .ZN(_16410_));
 MUX2_X1 _26134_ (.A(_01225_),
    .B(_16410_),
    .S(_16040_),
    .Z(_01074_));
 NAND4_X1 _26135_ (.A1(_16268_),
    .A2(_16221_),
    .A3(_16171_),
    .A4(_16270_),
    .ZN(_16411_));
 NAND2_X1 _26136_ (.A1(_16262_),
    .A2(_16411_),
    .ZN(_16412_));
 NOR2_X1 _26137_ (.A1(_16314_),
    .A2(_16283_),
    .ZN(_16413_));
 INV_X1 _26138_ (.A(_16413_),
    .ZN(_16414_));
 AOI211_X1 _26139_ (.A(_16254_),
    .B(_16412_),
    .C1(_16258_),
    .C2(_16414_),
    .ZN(_16415_));
 BUF_X2 _26140_ (.A(_16286_),
    .Z(_16416_));
 NAND2_X1 _26141_ (.A1(_16416_),
    .A2(_16317_),
    .ZN(_16417_));
 INV_X1 _26142_ (.A(_16286_),
    .ZN(_16418_));
 INV_X1 _26143_ (.A(_16318_),
    .ZN(_16419_));
 OAI21_X1 _26144_ (.A(_16417_),
    .B1(_16418_),
    .B2(_16419_),
    .ZN(_16420_));
 INV_X1 _26145_ (.A(_16197_),
    .ZN(_16421_));
 AOI211_X1 _26146_ (.A(_10986_),
    .B(_16418_),
    .C1(_16289_),
    .C2(_16421_),
    .ZN(_16422_));
 AOI211_X1 _26147_ (.A(_16420_),
    .B(_16422_),
    .C1(_16257_),
    .C2(_16416_),
    .ZN(_16423_));
 BUF_X2 _26148_ (.A(_16175_),
    .Z(_16424_));
 NAND3_X1 _26149_ (.A1(_16308_),
    .A2(_16424_),
    .A3(_16269_),
    .ZN(_16425_));
 BUF_X2 _26150_ (.A(_16223_),
    .Z(_16426_));
 AND2_X1 _26151_ (.A1(_16264_),
    .A2(_16426_),
    .ZN(_16427_));
 INV_X1 _26152_ (.A(_16427_),
    .ZN(_16428_));
 NAND2_X1 _26153_ (.A1(_16264_),
    .A2(_16302_),
    .ZN(_16429_));
 BUF_X2 _26154_ (.A(_16310_),
    .Z(_16430_));
 NAND2_X1 _26155_ (.A1(_16264_),
    .A2(_16430_),
    .ZN(_16431_));
 AND4_X1 _26156_ (.A1(_16425_),
    .A2(_16428_),
    .A3(_16429_),
    .A4(_16431_),
    .ZN(_16432_));
 NAND2_X1 _26157_ (.A1(_16281_),
    .A2(_16430_),
    .ZN(_16433_));
 CLKBUF_X2 _26158_ (.A(_16312_),
    .Z(_16434_));
 NAND2_X1 _26159_ (.A1(_16281_),
    .A2(_16434_),
    .ZN(_16435_));
 NAND2_X1 _26160_ (.A1(_16433_),
    .A2(_16435_),
    .ZN(_16436_));
 AND2_X1 _26161_ (.A1(_16281_),
    .A2(_16183_),
    .ZN(_16437_));
 AND2_X1 _26162_ (.A1(_16280_),
    .A2(_16344_),
    .ZN(_16438_));
 AND3_X1 _26163_ (.A1(_16306_),
    .A2(_16225_),
    .A3(_16268_),
    .ZN(_16439_));
 NOR4_X1 _26164_ (.A1(_16436_),
    .A2(_16437_),
    .A3(_16438_),
    .A4(_16439_),
    .ZN(_16440_));
 AND4_X1 _26165_ (.A1(_16415_),
    .A2(_16423_),
    .A3(_16432_),
    .A4(_16440_),
    .ZN(_16441_));
 AND2_X1 _26166_ (.A1(_16177_),
    .A2(_16211_),
    .ZN(_16442_));
 INV_X1 _26167_ (.A(_16442_),
    .ZN(_16443_));
 AND2_X1 _26168_ (.A1(_16177_),
    .A2(_16206_),
    .ZN(_16444_));
 INV_X1 _26169_ (.A(_16444_),
    .ZN(_16445_));
 NAND3_X1 _26170_ (.A1(_16377_),
    .A2(_16175_),
    .A3(_16176_),
    .ZN(_16446_));
 AND2_X1 _26171_ (.A1(_16189_),
    .A2(_16162_),
    .ZN(_16447_));
 NAND2_X1 _26172_ (.A1(_16178_),
    .A2(_16447_),
    .ZN(_16448_));
 AND4_X1 _26173_ (.A1(_16443_),
    .A2(_16445_),
    .A3(_16446_),
    .A4(_16448_),
    .ZN(_16449_));
 BUF_X2 _26174_ (.A(_16199_),
    .Z(_16450_));
 NAND2_X1 _26175_ (.A1(_16450_),
    .A2(_16426_),
    .ZN(_16451_));
 NAND2_X1 _26176_ (.A1(_16216_),
    .A2(_16190_),
    .ZN(_16452_));
 INV_X1 _26177_ (.A(_16452_),
    .ZN(_16453_));
 OAI21_X1 _26178_ (.A(_16450_),
    .B1(_16453_),
    .B2(_16183_),
    .ZN(_16454_));
 AND4_X1 _26179_ (.A1(_16208_),
    .A2(_16449_),
    .A3(_16451_),
    .A4(_16454_),
    .ZN(_16455_));
 OAI21_X1 _26180_ (.A(_16219_),
    .B1(_16453_),
    .B2(_16290_),
    .ZN(_16456_));
 CLKBUF_X2 _26181_ (.A(_16237_),
    .Z(_16457_));
 AOI21_X1 _26182_ (.A(_16243_),
    .B1(_16399_),
    .B2(_16457_),
    .ZN(_16458_));
 INV_X1 _26183_ (.A(_16245_),
    .ZN(_16459_));
 AND3_X1 _26184_ (.A1(_16237_),
    .A2(_16164_),
    .A3(_16167_),
    .ZN(_16460_));
 INV_X1 _26185_ (.A(_16460_),
    .ZN(_16461_));
 NAND2_X1 _26186_ (.A1(_16434_),
    .A2(_16237_),
    .ZN(_16462_));
 OAI211_X1 _26187_ (.A(_16237_),
    .B(_16426_),
    .C1(_16239_),
    .C2(_16276_),
    .ZN(_16463_));
 AND4_X1 _26188_ (.A1(_16459_),
    .A2(_16461_),
    .A3(_16462_),
    .A4(_16463_),
    .ZN(_16464_));
 AND4_X1 _26189_ (.A1(_16455_),
    .A2(_16456_),
    .A3(_16458_),
    .A4(_16464_),
    .ZN(_16465_));
 NOR2_X1 _26190_ (.A1(_16379_),
    .A2(_16452_),
    .ZN(_16466_));
 INV_X1 _26191_ (.A(_16466_),
    .ZN(_16467_));
 NAND4_X1 _26192_ (.A1(_16367_),
    .A2(_10987_),
    .A3(_16221_),
    .A4(_16270_),
    .ZN(_16468_));
 OAI21_X1 _26193_ (.A(_16371_),
    .B1(_16430_),
    .B2(_16207_),
    .ZN(_16469_));
 OAI211_X1 _26194_ (.A(_16371_),
    .B(_16426_),
    .C1(_16164_),
    .C2(_16171_),
    .ZN(_16470_));
 AND4_X1 _26195_ (.A1(_16467_),
    .A2(_16468_),
    .A3(_16469_),
    .A4(_16470_),
    .ZN(_16471_));
 INV_X1 _26196_ (.A(_16360_),
    .ZN(_16472_));
 NOR2_X1 _26197_ (.A1(_16472_),
    .A2(_16242_),
    .ZN(_16473_));
 INV_X1 _26198_ (.A(_16353_),
    .ZN(_16474_));
 INV_X1 _26199_ (.A(_16206_),
    .ZN(_16475_));
 OAI21_X1 _26200_ (.A(_16474_),
    .B1(_16472_),
    .B2(_16475_),
    .ZN(_16476_));
 BUF_X2 _26201_ (.A(_16360_),
    .Z(_16477_));
 AOI211_X1 _26202_ (.A(_16473_),
    .B(_16476_),
    .C1(_16477_),
    .C2(_16447_),
    .ZN(_16478_));
 AND2_X1 _26203_ (.A1(_16381_),
    .A2(_16310_),
    .ZN(_16479_));
 INV_X1 _26204_ (.A(_16479_),
    .ZN(_16480_));
 OAI21_X1 _26205_ (.A(_16381_),
    .B1(_16357_),
    .B2(_16299_),
    .ZN(_16481_));
 NAND3_X1 _26206_ (.A1(_16315_),
    .A2(_16175_),
    .A3(_16367_),
    .ZN(_16482_));
 BUF_X2 _26207_ (.A(_16224_),
    .Z(_16483_));
 OAI211_X1 _26208_ (.A(_16175_),
    .B(_16367_),
    .C1(_16275_),
    .C2(_16483_),
    .ZN(_16484_));
 AND4_X1 _26209_ (.A1(_16480_),
    .A2(_16481_),
    .A3(_16482_),
    .A4(_16484_),
    .ZN(_16485_));
 AND2_X1 _26210_ (.A1(_16182_),
    .A2(_10986_),
    .ZN(_16486_));
 NAND2_X1 _26211_ (.A1(_16390_),
    .A2(_16486_),
    .ZN(_16487_));
 NAND4_X1 _26212_ (.A1(_16190_),
    .A2(_16367_),
    .A3(_16236_),
    .A4(_16186_),
    .ZN(_16488_));
 NAND2_X1 _26213_ (.A1(_16487_),
    .A2(_16488_),
    .ZN(_16489_));
 AND2_X1 _26214_ (.A1(_16390_),
    .A2(_16223_),
    .ZN(_16490_));
 AOI221_X4 _26215_ (.A(_16489_),
    .B1(_16490_),
    .B2(_16187_),
    .C1(_16396_),
    .C2(_16414_),
    .ZN(_16491_));
 AND4_X1 _26216_ (.A1(_16471_),
    .A2(_16478_),
    .A3(_16485_),
    .A4(_16491_),
    .ZN(_16492_));
 BUF_X2 _26217_ (.A(_16305_),
    .Z(_16493_));
 OAI21_X1 _26218_ (.A(_16493_),
    .B1(_16220_),
    .B2(_16486_),
    .ZN(_16494_));
 NAND2_X1 _26219_ (.A1(_16354_),
    .A2(_16296_),
    .ZN(_16495_));
 AND2_X1 _26220_ (.A1(_16312_),
    .A2(_16339_),
    .ZN(_16496_));
 AND2_X1 _26221_ (.A1(_16354_),
    .A2(_16339_),
    .ZN(_16497_));
 AND2_X1 _26222_ (.A1(_16302_),
    .A2(_16339_),
    .ZN(_16498_));
 AND2_X1 _26223_ (.A1(_16339_),
    .A2(_16227_),
    .ZN(_16499_));
 NOR4_X1 _26224_ (.A1(_16496_),
    .A2(_16497_),
    .A3(_16498_),
    .A4(_16499_),
    .ZN(_16500_));
 OAI211_X1 _26225_ (.A(_16296_),
    .B(_16230_),
    .C1(_16239_),
    .C2(_16276_),
    .ZN(_16501_));
 OAI21_X1 _26226_ (.A(_16295_),
    .B1(_16275_),
    .B2(_16224_),
    .ZN(_16502_));
 AND4_X1 _26227_ (.A1(_16495_),
    .A2(_16500_),
    .A3(_16501_),
    .A4(_16502_),
    .ZN(_16503_));
 AND2_X1 _26228_ (.A1(_16312_),
    .A2(_16322_),
    .ZN(_16504_));
 AND2_X1 _26229_ (.A1(_16228_),
    .A2(_16322_),
    .ZN(_16505_));
 AND2_X1 _26230_ (.A1(_16322_),
    .A2(_16224_),
    .ZN(_16506_));
 NOR3_X1 _26231_ (.A1(_16504_),
    .A2(_16505_),
    .A3(_16506_),
    .ZN(_16507_));
 BUF_X2 _26232_ (.A(_16322_),
    .Z(_16508_));
 OAI21_X1 _26233_ (.A(_16508_),
    .B1(_16397_),
    .B2(_16299_),
    .ZN(_16509_));
 BUF_X2 _26234_ (.A(_16190_),
    .Z(_16510_));
 NAND4_X1 _26235_ (.A1(_16510_),
    .A2(_10987_),
    .A3(_16327_),
    .A4(_16270_),
    .ZN(_16511_));
 AND3_X1 _26236_ (.A1(_16507_),
    .A2(_16509_),
    .A3(_16511_),
    .ZN(_16512_));
 AND2_X1 _26237_ (.A1(_16305_),
    .A2(_16315_),
    .ZN(_16513_));
 AND2_X1 _26238_ (.A1(_16305_),
    .A2(_16227_),
    .ZN(_16514_));
 AOI221_X4 _26239_ (.A(_16513_),
    .B1(_16305_),
    .B2(_16224_),
    .C1(_10986_),
    .C2(_16514_),
    .ZN(_16515_));
 AND4_X1 _26240_ (.A1(_16494_),
    .A2(_16503_),
    .A3(_16512_),
    .A4(_16515_),
    .ZN(_16516_));
 NAND4_X1 _26241_ (.A1(_16441_),
    .A2(_16465_),
    .A3(_16492_),
    .A4(_16516_),
    .ZN(_16517_));
 NOR2_X1 _26242_ (.A1(_16517_),
    .A2(_16406_),
    .ZN(_16518_));
 XOR2_X1 _26243_ (.A(_01016_),
    .B(_01015_),
    .Z(_16519_));
 XNOR2_X1 _26244_ (.A(_16518_),
    .B(_16519_),
    .ZN(_16520_));
 MUX2_X1 _26245_ (.A(_01226_),
    .B(_16520_),
    .S(_16040_),
    .Z(_01075_));
 AND2_X1 _26246_ (.A1(_16207_),
    .A2(_16348_),
    .ZN(_16521_));
 INV_X1 _26247_ (.A(_16170_),
    .ZN(_16522_));
 AND3_X1 _26248_ (.A1(_16290_),
    .A2(_16348_),
    .A3(_16522_),
    .ZN(_16523_));
 AND4_X1 _26249_ (.A1(_10986_),
    .A2(_16327_),
    .A3(_16223_),
    .A4(_16236_),
    .ZN(_16524_));
 OR4_X1 _26250_ (.A1(_16521_),
    .A2(_16523_),
    .A3(_16498_),
    .A4(_16524_),
    .ZN(_16525_));
 AND2_X1 _26251_ (.A1(_16296_),
    .A2(_16197_),
    .ZN(_16526_));
 NOR2_X1 _26252_ (.A1(_16234_),
    .A2(_16170_),
    .ZN(_16527_));
 AND2_X1 _26253_ (.A1(_16527_),
    .A2(_16295_),
    .ZN(_16528_));
 AOI21_X1 _26254_ (.A(_16335_),
    .B1(_16334_),
    .B2(_16284_),
    .ZN(_16529_));
 NOR4_X1 _26255_ (.A1(_16525_),
    .A2(_16526_),
    .A3(_16528_),
    .A4(_16529_),
    .ZN(_16530_));
 NAND2_X1 _26256_ (.A1(_16493_),
    .A2(_16197_),
    .ZN(_16531_));
 NAND2_X1 _26257_ (.A1(_16493_),
    .A2(_16344_),
    .ZN(_16532_));
 NAND2_X1 _26258_ (.A1(_16493_),
    .A2(_16183_),
    .ZN(_16533_));
 AND3_X1 _26259_ (.A1(_16531_),
    .A2(_16532_),
    .A3(_16533_),
    .ZN(_16534_));
 NAND3_X1 _26260_ (.A1(_16483_),
    .A2(_16424_),
    .A3(_16327_),
    .ZN(_16535_));
 INV_X1 _26261_ (.A(_16514_),
    .ZN(_16536_));
 OAI21_X1 _26262_ (.A(_16493_),
    .B1(_16315_),
    .B2(_16283_),
    .ZN(_16537_));
 NAND4_X1 _26263_ (.A1(_16534_),
    .A2(_16535_),
    .A3(_16536_),
    .A4(_16537_),
    .ZN(_16538_));
 OAI211_X1 _26264_ (.A(_16508_),
    .B(_16510_),
    .C1(_16164_),
    .C2(_16186_),
    .ZN(_16539_));
 INV_X1 _26265_ (.A(_16322_),
    .ZN(_16540_));
 OAI21_X1 _26266_ (.A(_16539_),
    .B1(_16540_),
    .B2(_16421_),
    .ZN(_16541_));
 NAND3_X1 _26267_ (.A1(_16508_),
    .A2(_16230_),
    .A3(_16187_),
    .ZN(_16542_));
 NAND2_X1 _26268_ (.A1(_16321_),
    .A2(_16542_),
    .ZN(_16543_));
 INV_X1 _26269_ (.A(_16308_),
    .ZN(_16544_));
 AOI21_X1 _26270_ (.A(_16540_),
    .B1(_16544_),
    .B2(_16298_),
    .ZN(_16545_));
 NOR4_X1 _26271_ (.A1(_16538_),
    .A2(_16541_),
    .A3(_16543_),
    .A4(_16545_),
    .ZN(_16546_));
 AND2_X1 _26272_ (.A1(_16250_),
    .A2(_16206_),
    .ZN(_16547_));
 INV_X1 _26273_ (.A(_16547_),
    .ZN(_16548_));
 NAND3_X1 _26274_ (.A1(_16430_),
    .A2(_16269_),
    .A3(_16270_),
    .ZN(_16549_));
 NAND2_X1 _26275_ (.A1(_16250_),
    .A2(_16277_),
    .ZN(_16550_));
 NAND3_X1 _26276_ (.A1(_16548_),
    .A2(_16549_),
    .A3(_16550_),
    .ZN(_16551_));
 NAND2_X1 _26277_ (.A1(_16264_),
    .A2(_16183_),
    .ZN(_16552_));
 NAND2_X1 _26278_ (.A1(_16264_),
    .A2(_16278_),
    .ZN(_16553_));
 NAND3_X1 _26279_ (.A1(_16434_),
    .A2(_16424_),
    .A3(_16269_),
    .ZN(_16554_));
 NAND4_X1 _26280_ (.A1(_16552_),
    .A2(_16431_),
    .A3(_16553_),
    .A4(_16554_),
    .ZN(_16555_));
 OAI21_X1 _26281_ (.A(_16221_),
    .B1(_10986_),
    .B2(_16276_),
    .ZN(_16556_));
 INV_X1 _26282_ (.A(_16556_),
    .ZN(_16557_));
 AND2_X1 _26283_ (.A1(_16258_),
    .A2(_16557_),
    .ZN(_16558_));
 NAND2_X1 _26284_ (.A1(_16258_),
    .A2(_16273_),
    .ZN(_16559_));
 NAND2_X1 _26285_ (.A1(_16258_),
    .A2(_16306_),
    .ZN(_16560_));
 NAND4_X1 _26286_ (.A1(_16269_),
    .A2(_10993_),
    .A3(_16510_),
    .A4(_16270_),
    .ZN(_16561_));
 NAND3_X1 _26287_ (.A1(_16559_),
    .A2(_16560_),
    .A3(_16561_),
    .ZN(_16562_));
 NOR4_X1 _26288_ (.A1(_16551_),
    .A2(_16555_),
    .A3(_16558_),
    .A4(_16562_),
    .ZN(_16563_));
 AOI211_X1 _26289_ (.A(_16260_),
    .B(_16418_),
    .C1(_10987_),
    .C2(_10993_),
    .ZN(_16564_));
 OAI21_X1 _26290_ (.A(_16281_),
    .B1(_16306_),
    .B2(_16197_),
    .ZN(_16565_));
 NAND2_X1 _26291_ (.A1(_16281_),
    .A2(_16315_),
    .ZN(_16566_));
 OAI211_X1 _26292_ (.A(_16565_),
    .B(_16566_),
    .C1(_16213_),
    .C2(_16282_),
    .ZN(_16567_));
 NAND2_X1 _26293_ (.A1(_16416_),
    .A2(_16483_),
    .ZN(_16568_));
 NAND3_X1 _26294_ (.A1(_16430_),
    .A2(_16268_),
    .A3(_16236_),
    .ZN(_16569_));
 NAND4_X1 _26295_ (.A1(_16269_),
    .A2(_16171_),
    .A3(_16230_),
    .A4(_16236_),
    .ZN(_16570_));
 NAND4_X1 _26296_ (.A1(_16568_),
    .A2(_16417_),
    .A3(_16569_),
    .A4(_16570_),
    .ZN(_16571_));
 NOR4_X1 _26297_ (.A1(_16564_),
    .A2(_16567_),
    .A3(_16291_),
    .A4(_16571_),
    .ZN(_16572_));
 NAND4_X1 _26298_ (.A1(_16530_),
    .A2(_16546_),
    .A3(_16563_),
    .A4(_16572_),
    .ZN(_16573_));
 NAND3_X1 _26299_ (.A1(_16434_),
    .A2(_16424_),
    .A3(_16176_),
    .ZN(_16574_));
 OAI21_X1 _26300_ (.A(_16178_),
    .B1(_16283_),
    .B2(_16244_),
    .ZN(_16575_));
 OAI21_X1 _26301_ (.A(_16180_),
    .B1(_16354_),
    .B2(_16397_),
    .ZN(_16576_));
 NAND3_X1 _26302_ (.A1(_16278_),
    .A2(_16175_),
    .A3(_16176_),
    .ZN(_16577_));
 AND4_X1 _26303_ (.A1(_16574_),
    .A2(_16575_),
    .A3(_16576_),
    .A4(_16577_),
    .ZN(_16578_));
 NAND3_X1 _26304_ (.A1(_16265_),
    .A2(_16187_),
    .A3(_16450_),
    .ZN(_16579_));
 AND2_X1 _26305_ (.A1(_16527_),
    .A2(_16199_),
    .ZN(_16580_));
 AND3_X1 _26306_ (.A1(_16199_),
    .A2(_16171_),
    .A3(_16167_),
    .ZN(_16581_));
 NOR2_X1 _26307_ (.A1(_16580_),
    .A2(_16581_),
    .ZN(_16582_));
 AND4_X1 _26308_ (.A1(_16201_),
    .A2(_16578_),
    .A3(_16579_),
    .A4(_16582_),
    .ZN(_16583_));
 NAND2_X1 _26309_ (.A1(_16172_),
    .A2(_16477_),
    .ZN(_16584_));
 OAI21_X1 _26310_ (.A(_16477_),
    .B1(_16317_),
    .B2(_16318_),
    .ZN(_16585_));
 OAI211_X1 _26311_ (.A(_16477_),
    .B(_16510_),
    .C1(_16164_),
    .C2(_16193_),
    .ZN(_16586_));
 NAND4_X1 _26312_ (.A1(_16584_),
    .A2(_16363_),
    .A3(_16585_),
    .A4(_16586_),
    .ZN(_16587_));
 NAND2_X1 _26313_ (.A1(_16400_),
    .A2(_16398_),
    .ZN(_16588_));
 AND2_X1 _26314_ (.A1(_16310_),
    .A2(_16396_),
    .ZN(_16589_));
 NOR4_X1 _26315_ (.A1(_16587_),
    .A2(_16393_),
    .A3(_16588_),
    .A4(_16589_),
    .ZN(_16590_));
 OAI21_X1 _26316_ (.A(_16375_),
    .B1(_16306_),
    .B2(_16308_),
    .ZN(_16591_));
 OAI21_X1 _26317_ (.A(_16385_),
    .B1(_16306_),
    .B2(_16397_),
    .ZN(_16592_));
 OAI21_X1 _26318_ (.A(_16385_),
    .B1(_16315_),
    .B2(_16331_),
    .ZN(_16593_));
 OAI21_X1 _26319_ (.A(_16375_),
    .B1(_16315_),
    .B2(_16228_),
    .ZN(_16594_));
 AND4_X1 _26320_ (.A1(_16591_),
    .A2(_16592_),
    .A3(_16593_),
    .A4(_16594_),
    .ZN(_16595_));
 OAI21_X1 _26321_ (.A(_16457_),
    .B1(_16244_),
    .B2(_16331_),
    .ZN(_16596_));
 NAND4_X1 _26322_ (.A1(_16457_),
    .A2(_16510_),
    .A3(_16216_),
    .A4(_16187_),
    .ZN(_16597_));
 OAI211_X1 _26323_ (.A(_16596_),
    .B(_16597_),
    .C1(_16238_),
    .C2(_16378_),
    .ZN(_16598_));
 NAND2_X1 _26324_ (.A1(_16219_),
    .A2(_16430_),
    .ZN(_16599_));
 NAND4_X1 _26325_ (.A1(_16225_),
    .A2(_16426_),
    .A3(_16193_),
    .A4(_16176_),
    .ZN(_16600_));
 INV_X1 _26326_ (.A(_16218_),
    .ZN(_16601_));
 OAI211_X1 _26327_ (.A(_16599_),
    .B(_16600_),
    .C1(_16334_),
    .C2(_16601_),
    .ZN(_16602_));
 NAND2_X1 _26328_ (.A1(_16219_),
    .A2(_16302_),
    .ZN(_16603_));
 OAI21_X1 _26329_ (.A(_16603_),
    .B1(_16601_),
    .B2(_16421_),
    .ZN(_16604_));
 AND2_X1 _26330_ (.A1(_16219_),
    .A2(_16557_),
    .ZN(_16605_));
 NOR4_X1 _26331_ (.A1(_16598_),
    .A2(_16602_),
    .A3(_16604_),
    .A4(_16605_),
    .ZN(_16606_));
 NAND4_X1 _26332_ (.A1(_16583_),
    .A2(_16590_),
    .A3(_16595_),
    .A4(_16606_),
    .ZN(_16607_));
 NOR2_X1 _26333_ (.A1(_16573_),
    .A2(_16607_),
    .ZN(_16608_));
 XOR2_X1 _26334_ (.A(_01018_),
    .B(_01017_),
    .Z(_16609_));
 XNOR2_X1 _26335_ (.A(_16608_),
    .B(_16609_),
    .ZN(_16610_));
 MUX2_X1 _26336_ (.A(_01227_),
    .B(_16610_),
    .S(_16040_),
    .Z(_01076_));
 AND2_X1 _26337_ (.A1(_16416_),
    .A2(_16318_),
    .ZN(_16611_));
 AND4_X1 _26338_ (.A1(_16165_),
    .A2(_16286_),
    .A3(_16522_),
    .A4(_16167_),
    .ZN(_16612_));
 AOI211_X1 _26339_ (.A(_16611_),
    .B(_16612_),
    .C1(_16228_),
    .C2(_16416_),
    .ZN(_16613_));
 NAND4_X1 _26340_ (.A1(_16269_),
    .A2(_10987_),
    .A3(_16236_),
    .A4(_16221_),
    .ZN(_16614_));
 OAI211_X1 _26341_ (.A(_16416_),
    .B(_16510_),
    .C1(_16239_),
    .C2(_10993_),
    .ZN(_16615_));
 NAND3_X1 _26342_ (.A1(_16613_),
    .A2(_16614_),
    .A3(_16615_),
    .ZN(_16616_));
 NOR3_X1 _26343_ (.A1(_16163_),
    .A2(_16188_),
    .A3(_17077_),
    .ZN(_16617_));
 NAND3_X1 _26344_ (.A1(_16493_),
    .A2(_16522_),
    .A3(_16617_),
    .ZN(_16618_));
 NAND2_X1 _26345_ (.A1(_16434_),
    .A2(_16450_),
    .ZN(_16619_));
 NAND2_X1 _26346_ (.A1(_16317_),
    .A2(_16450_),
    .ZN(_16620_));
 NAND3_X1 _26347_ (.A1(_16618_),
    .A2(_16619_),
    .A3(_16620_),
    .ZN(_16621_));
 INV_X1 _26348_ (.A(_16486_),
    .ZN(_16622_));
 AOI21_X1 _26349_ (.A(_16204_),
    .B1(_16195_),
    .B2(_16622_),
    .ZN(_16623_));
 AND2_X1 _26350_ (.A1(_16167_),
    .A2(_16162_),
    .ZN(_16624_));
 INV_X1 _26351_ (.A(_16624_),
    .ZN(_16625_));
 AOI21_X1 _26352_ (.A(_16391_),
    .B1(_16195_),
    .B2(_16625_),
    .ZN(_16626_));
 NOR4_X1 _26353_ (.A1(_16616_),
    .A2(_16621_),
    .A3(_16623_),
    .A4(_16626_),
    .ZN(_16627_));
 NAND2_X1 _26354_ (.A1(_16180_),
    .A2(_16302_),
    .ZN(_16628_));
 AOI22_X1 _26355_ (.A1(_16180_),
    .A2(_16483_),
    .B1(_16273_),
    .B2(_16508_),
    .ZN(_16629_));
 NAND2_X1 _26356_ (.A1(_16385_),
    .A2(_16207_),
    .ZN(_16630_));
 NAND2_X1 _26357_ (.A1(_16483_),
    .A2(_16457_),
    .ZN(_16631_));
 AND4_X1 _26358_ (.A1(_16628_),
    .A2(_16629_),
    .A3(_16630_),
    .A4(_16631_),
    .ZN(_16632_));
 AOI21_X1 _26359_ (.A(_16346_),
    .B1(_16284_),
    .B2(_16300_),
    .ZN(_16633_));
 AND2_X1 _26360_ (.A1(_16360_),
    .A2(_16318_),
    .ZN(_16634_));
 AND2_X1 _26361_ (.A1(_16397_),
    .A2(_16322_),
    .ZN(_16635_));
 NOR4_X1 _26362_ (.A1(_16633_),
    .A2(_16634_),
    .A3(_16393_),
    .A4(_16635_),
    .ZN(_16636_));
 OAI21_X1 _26363_ (.A(_16399_),
    .B1(_16264_),
    .B2(_16218_),
    .ZN(_16637_));
 NAND2_X1 _26364_ (.A1(_16318_),
    .A2(_16218_),
    .ZN(_16638_));
 NAND3_X1 _26365_ (.A1(_16617_),
    .A2(_16522_),
    .A3(_16237_),
    .ZN(_16639_));
 AND4_X1 _26366_ (.A1(_16559_),
    .A2(_16637_),
    .A3(_16638_),
    .A4(_16639_),
    .ZN(_16640_));
 NAND2_X1 _26367_ (.A1(_16344_),
    .A2(_16218_),
    .ZN(_16641_));
 NAND4_X1 _26368_ (.A1(_16228_),
    .A2(_10986_),
    .A3(_16225_),
    .A4(_16268_),
    .ZN(_16642_));
 NAND2_X1 _26369_ (.A1(_16308_),
    .A2(_16296_),
    .ZN(_16643_));
 AND4_X1 _26370_ (.A1(_16641_),
    .A2(_16642_),
    .A3(_16643_),
    .A4(_16398_),
    .ZN(_16644_));
 AND4_X1 _26371_ (.A1(_16632_),
    .A2(_16636_),
    .A3(_16640_),
    .A4(_16644_),
    .ZN(_16645_));
 AND2_X1 _26372_ (.A1(_16302_),
    .A2(_16295_),
    .ZN(_16646_));
 AND2_X1 _26373_ (.A1(_16223_),
    .A2(_16162_),
    .ZN(_16647_));
 AND2_X1 _26374_ (.A1(_16371_),
    .A2(_16647_),
    .ZN(_16648_));
 AND2_X1 _26375_ (.A1(_16322_),
    .A2(_16377_),
    .ZN(_16649_));
 NOR4_X1 _26376_ (.A1(_16479_),
    .A2(_16646_),
    .A3(_16648_),
    .A4(_16649_),
    .ZN(_16650_));
 AOI221_X4 _26377_ (.A(_16382_),
    .B1(_16183_),
    .B2(_16348_),
    .C1(_16278_),
    .C2(_16508_),
    .ZN(_16651_));
 NAND2_X1 _26378_ (.A1(_16381_),
    .A2(_16426_),
    .ZN(_16652_));
 NAND2_X1 _26379_ (.A1(_16178_),
    .A2(_16290_),
    .ZN(_16653_));
 AND4_X1 _26380_ (.A1(_16552_),
    .A2(_16428_),
    .A3(_16652_),
    .A4(_16653_),
    .ZN(_16654_));
 NAND2_X1 _26381_ (.A1(_16381_),
    .A2(_16399_),
    .ZN(_16655_));
 AOI22_X1 _26382_ (.A1(_16228_),
    .A2(_16360_),
    .B1(_16430_),
    .B2(_16322_),
    .ZN(_16656_));
 AND3_X1 _26383_ (.A1(_16548_),
    .A2(_16655_),
    .A3(_16656_),
    .ZN(_16657_));
 AND4_X1 _26384_ (.A1(_16650_),
    .A2(_16651_),
    .A3(_16654_),
    .A4(_16657_),
    .ZN(_16658_));
 AND2_X1 _26385_ (.A1(_16295_),
    .A2(_16483_),
    .ZN(_16659_));
 NOR4_X1 _26386_ (.A1(_16473_),
    .A2(_16521_),
    .A3(_16340_),
    .A4(_16659_),
    .ZN(_16660_));
 AOI22_X1 _26387_ (.A1(_16325_),
    .A2(_10993_),
    .B1(_16258_),
    .B2(_16557_),
    .ZN(_16661_));
 AND4_X1 _26388_ (.A1(_16467_),
    .A2(_16660_),
    .A3(_16495_),
    .A4(_16661_),
    .ZN(_16662_));
 NAND4_X1 _26389_ (.A1(_16627_),
    .A2(_16645_),
    .A3(_16658_),
    .A4(_16662_),
    .ZN(_16663_));
 INV_X1 _26390_ (.A(_16313_),
    .ZN(_16664_));
 OAI21_X1 _26391_ (.A(_16296_),
    .B1(_16344_),
    .B2(_16228_),
    .ZN(_16665_));
 AND3_X1 _26392_ (.A1(_16664_),
    .A2(_16536_),
    .A3(_16665_),
    .ZN(_16666_));
 NAND2_X1 _26393_ (.A1(_16477_),
    .A2(_16257_),
    .ZN(_16667_));
 OAI21_X1 _26394_ (.A(_16375_),
    .B1(_16283_),
    .B2(_16290_),
    .ZN(_16668_));
 AND4_X1 _26395_ (.A1(_16342_),
    .A2(_16666_),
    .A3(_16667_),
    .A4(_16668_),
    .ZN(_16669_));
 AND2_X1 _26396_ (.A1(_16280_),
    .A2(_16357_),
    .ZN(_16670_));
 NOR2_X1 _26397_ (.A1(_16670_),
    .A2(_16274_),
    .ZN(_16671_));
 INV_X1 _26398_ (.A(_16263_),
    .ZN(_16672_));
 OR2_X1 _26399_ (.A1(_16413_),
    .A2(_16672_),
    .ZN(_16673_));
 AND2_X1 _26400_ (.A1(_16434_),
    .A2(_16296_),
    .ZN(_16674_));
 AND2_X1 _26401_ (.A1(_16357_),
    .A2(_16339_),
    .ZN(_16675_));
 NOR2_X1 _26402_ (.A1(_16674_),
    .A2(_16675_),
    .ZN(_16676_));
 NAND2_X1 _26403_ (.A1(_16483_),
    .A2(_16450_),
    .ZN(_16677_));
 AND2_X1 _26404_ (.A1(_16566_),
    .A2(_16677_),
    .ZN(_01332_));
 AND4_X1 _26405_ (.A1(_16671_),
    .A2(_16673_),
    .A3(_16676_),
    .A4(_01332_),
    .ZN(_01333_));
 INV_X1 _26406_ (.A(_16213_),
    .ZN(_01334_));
 AOI22_X1 _26407_ (.A1(_01334_),
    .A2(_16258_),
    .B1(_16180_),
    .B2(_16172_),
    .ZN(_01335_));
 INV_X1 _26408_ (.A(_16306_),
    .ZN(_01336_));
 OAI21_X1 _26409_ (.A(_16532_),
    .B1(_01336_),
    .B2(_16472_),
    .ZN(_01337_));
 AND2_X1 _26410_ (.A1(_16430_),
    .A2(_16296_),
    .ZN(_01338_));
 NOR4_X1 _26411_ (.A1(_01337_),
    .A2(_16437_),
    .A3(_01338_),
    .A4(_16505_),
    .ZN(_01339_));
 NAND4_X1 _26412_ (.A1(_16669_),
    .A2(_01333_),
    .A3(_01335_),
    .A4(_01339_),
    .ZN(_01340_));
 NOR2_X1 _26413_ (.A1(_16663_),
    .A2(_01340_),
    .ZN(_01341_));
 XOR2_X1 _26414_ (.A(_01020_),
    .B(_01019_),
    .Z(_01342_));
 XNOR2_X1 _26415_ (.A(_01341_),
    .B(_01342_),
    .ZN(_01343_));
 MUX2_X1 _26416_ (.A(_01228_),
    .B(_01343_),
    .S(_16040_),
    .Z(_01077_));
 AOI211_X1 _26417_ (.A(_16193_),
    .B(_16601_),
    .C1(_16260_),
    .C2(_16289_),
    .ZN(_01344_));
 NOR3_X1 _26418_ (.A1(_16601_),
    .A2(_16171_),
    .A3(_16168_),
    .ZN(_01345_));
 AND2_X1 _26419_ (.A1(_16218_),
    .A2(_16278_),
    .ZN(_01346_));
 OR3_X1 _26420_ (.A1(_01345_),
    .A2(_16229_),
    .A3(_01346_),
    .ZN(_01347_));
 AND2_X1 _26421_ (.A1(_16228_),
    .A2(_16237_),
    .ZN(_01348_));
 OR2_X1 _26422_ (.A1(_16460_),
    .A2(_01348_),
    .ZN(_01349_));
 AND2_X1 _26423_ (.A1(_16261_),
    .A2(_16457_),
    .ZN(_01350_));
 NOR4_X1 _26424_ (.A1(_01344_),
    .A2(_01347_),
    .A3(_01349_),
    .A4(_01350_),
    .ZN(_01351_));
 OAI21_X1 _26425_ (.A(_16477_),
    .B1(_16283_),
    .B2(_16434_),
    .ZN(_01352_));
 NAND3_X1 _26426_ (.A1(_16477_),
    .A2(_16290_),
    .A3(_16522_),
    .ZN(_01353_));
 OAI211_X1 _26427_ (.A(_16477_),
    .B(_16426_),
    .C1(_16239_),
    .C2(_16276_),
    .ZN(_01354_));
 NAND4_X1 _26428_ (.A1(_16356_),
    .A2(_01352_),
    .A3(_01353_),
    .A4(_01354_),
    .ZN(_01355_));
 AND2_X1 _26429_ (.A1(_16315_),
    .A2(_16396_),
    .ZN(_01356_));
 OR2_X1 _26430_ (.A1(_16589_),
    .A2(_01356_),
    .ZN(_01357_));
 AOI21_X1 _26431_ (.A(_16391_),
    .B1(_16260_),
    .B2(_16300_),
    .ZN(_01358_));
 NOR4_X1 _26432_ (.A1(_01355_),
    .A2(_01357_),
    .A3(_16490_),
    .A4(_01358_),
    .ZN(_01359_));
 INV_X1 _26433_ (.A(_16383_),
    .ZN(_01360_));
 OAI21_X1 _26434_ (.A(_16385_),
    .B1(_16306_),
    .B2(_16197_),
    .ZN(_01361_));
 AND2_X1 _26435_ (.A1(_01360_),
    .A2(_01361_),
    .ZN(_01362_));
 NAND2_X1 _26436_ (.A1(_16354_),
    .A2(_16375_),
    .ZN(_01363_));
 NAND3_X1 _26437_ (.A1(_16397_),
    .A2(_16270_),
    .A3(_16367_),
    .ZN(_01364_));
 AND3_X1 _26438_ (.A1(_16376_),
    .A2(_01363_),
    .A3(_01364_),
    .ZN(_01365_));
 OAI21_X1 _26439_ (.A(_16385_),
    .B1(_16317_),
    .B2(_16207_),
    .ZN(_01366_));
 AND4_X1 _26440_ (.A1(_16469_),
    .A2(_01362_),
    .A3(_01365_),
    .A4(_01366_),
    .ZN(_01367_));
 OAI21_X1 _26441_ (.A(_16180_),
    .B1(_16302_),
    .B2(_16357_),
    .ZN(_01368_));
 OAI21_X1 _26442_ (.A(_16180_),
    .B1(_16317_),
    .B2(_16483_),
    .ZN(_01369_));
 NAND2_X1 _26443_ (.A1(_16180_),
    .A2(_16397_),
    .ZN(_01370_));
 NAND2_X1 _26444_ (.A1(_16178_),
    .A2(_16283_),
    .ZN(_01371_));
 NAND4_X1 _26445_ (.A1(_01368_),
    .A2(_01369_),
    .A3(_01370_),
    .A4(_01371_),
    .ZN(_01372_));
 INV_X1 _26446_ (.A(_16244_),
    .ZN(_01373_));
 OAI22_X1 _26447_ (.A1(_01373_),
    .A2(_16204_),
    .B1(_16451_),
    .B2(_16171_),
    .ZN(_01374_));
 INV_X1 _26448_ (.A(_16343_),
    .ZN(_01375_));
 AOI21_X1 _26449_ (.A(_16204_),
    .B1(_01375_),
    .B2(_16203_),
    .ZN(_01376_));
 AND3_X1 _26450_ (.A1(_16450_),
    .A2(_16510_),
    .A3(_16186_),
    .ZN(_01377_));
 NOR4_X1 _26451_ (.A1(_01372_),
    .A2(_01374_),
    .A3(_01376_),
    .A4(_01377_),
    .ZN(_01378_));
 NAND4_X1 _26452_ (.A1(_01351_),
    .A2(_01359_),
    .A3(_01367_),
    .A4(_01378_),
    .ZN(_01379_));
 AND3_X1 _26453_ (.A1(_16308_),
    .A2(_16225_),
    .A3(_16268_),
    .ZN(_01380_));
 OR3_X1 _26454_ (.A1(_16438_),
    .A2(_16670_),
    .A3(_01380_),
    .ZN(_01381_));
 AOI21_X1 _26455_ (.A(_16418_),
    .B1(_01336_),
    .B2(_16544_),
    .ZN(_01382_));
 AOI21_X1 _26456_ (.A(_16418_),
    .B1(_16413_),
    .B2(_16419_),
    .ZN(_01383_));
 NOR4_X1 _26457_ (.A1(_01381_),
    .A2(_16285_),
    .A3(_01382_),
    .A4(_01383_),
    .ZN(_01384_));
 AND2_X1 _26458_ (.A1(_16305_),
    .A2(_16354_),
    .ZN(_01385_));
 INV_X1 _26459_ (.A(_01385_),
    .ZN(_01386_));
 OAI21_X1 _26460_ (.A(_16493_),
    .B1(_16308_),
    .B2(_16377_),
    .ZN(_01387_));
 OAI211_X1 _26461_ (.A(_16493_),
    .B(_16230_),
    .C1(_10987_),
    .C2(_10993_),
    .ZN(_01388_));
 NAND4_X1 _26462_ (.A1(_01386_),
    .A2(_16536_),
    .A3(_01387_),
    .A4(_01388_),
    .ZN(_01389_));
 AND2_X1 _26463_ (.A1(_16447_),
    .A2(_16508_),
    .ZN(_01390_));
 NOR4_X1 _26464_ (.A1(_01389_),
    .A2(_16543_),
    .A3(_16649_),
    .A4(_01390_),
    .ZN(_01391_));
 OAI21_X1 _26465_ (.A(_16264_),
    .B1(_16354_),
    .B2(_16397_),
    .ZN(_01392_));
 NAND2_X1 _26466_ (.A1(_16264_),
    .A2(_16527_),
    .ZN(_01393_));
 OAI211_X1 _26467_ (.A(_01392_),
    .B(_01393_),
    .C1(_16475_),
    .C2(_16672_),
    .ZN(_01394_));
 NOR4_X1 _26468_ (.A1(_16256_),
    .A2(_01394_),
    .A3(_16412_),
    .A4(_16547_),
    .ZN(_01395_));
 NAND2_X1 _26469_ (.A1(_16348_),
    .A2(_16426_),
    .ZN(_01396_));
 OAI211_X1 _26470_ (.A(_16342_),
    .B(_01396_),
    .C1(_16284_),
    .C2(_16346_),
    .ZN(_01397_));
 NAND2_X1 _26471_ (.A1(_16344_),
    .A2(_16296_),
    .ZN(_01398_));
 NAND4_X1 _26472_ (.A1(_16225_),
    .A2(_10993_),
    .A3(_16327_),
    .A4(_16221_),
    .ZN(_01399_));
 NAND4_X1 _26473_ (.A1(_16510_),
    .A2(_16225_),
    .A3(_10987_),
    .A4(_16327_),
    .ZN(_01400_));
 NAND3_X1 _26474_ (.A1(_01398_),
    .A2(_01399_),
    .A3(_01400_),
    .ZN(_01401_));
 NOR4_X1 _26475_ (.A1(_01397_),
    .A2(_16332_),
    .A3(_01338_),
    .A4(_01401_),
    .ZN(_01402_));
 NAND4_X1 _26476_ (.A1(_01384_),
    .A2(_01391_),
    .A3(_01395_),
    .A4(_01402_),
    .ZN(_01403_));
 NOR2_X1 _26477_ (.A1(_01379_),
    .A2(_01403_),
    .ZN(_01404_));
 XOR2_X1 _26478_ (.A(_01022_),
    .B(_01021_),
    .Z(_01405_));
 XNOR2_X1 _26479_ (.A(_01404_),
    .B(_01405_),
    .ZN(_01406_));
 MUX2_X1 _26480_ (.A(_01229_),
    .B(_01406_),
    .S(_16040_),
    .Z(_01078_));
 OAI21_X1 _26481_ (.A(_16219_),
    .B1(_16647_),
    .B2(_16230_),
    .ZN(_01407_));
 AOI21_X1 _26482_ (.A(_01376_),
    .B1(_16450_),
    .B2(_16453_),
    .ZN(_01408_));
 AND2_X1 _26483_ (.A1(_16178_),
    .A2(_16244_),
    .ZN(_01409_));
 AOI211_X1 _26484_ (.A(_16444_),
    .B(_01409_),
    .C1(_01334_),
    .C2(_16178_),
    .ZN(_01410_));
 OAI221_X1 _26485_ (.A(_16450_),
    .B1(_16239_),
    .B2(_17075_),
    .C1(_16230_),
    .C2(_16426_),
    .ZN(_01411_));
 AND2_X1 _26486_ (.A1(_16617_),
    .A2(_16522_),
    .ZN(_01412_));
 OAI21_X1 _26487_ (.A(_16180_),
    .B1(_01412_),
    .B2(_16397_),
    .ZN(_01413_));
 AND4_X1 _26488_ (.A1(_01408_),
    .A2(_01410_),
    .A3(_01411_),
    .A4(_01413_),
    .ZN(_01414_));
 OAI21_X1 _26489_ (.A(_16219_),
    .B1(_16453_),
    .B2(_16557_),
    .ZN(_01415_));
 AND2_X1 _26490_ (.A1(_16308_),
    .A2(_16457_),
    .ZN(_01416_));
 AND2_X1 _26491_ (.A1(_16434_),
    .A2(_16457_),
    .ZN(_01417_));
 AND2_X1 _26492_ (.A1(_16278_),
    .A2(_16237_),
    .ZN(_01418_));
 NOR4_X1 _26493_ (.A1(_01416_),
    .A2(_01417_),
    .A3(_01418_),
    .A4(_01348_),
    .ZN(_01419_));
 AND4_X1 _26494_ (.A1(_01407_),
    .A2(_01414_),
    .A3(_01415_),
    .A4(_01419_),
    .ZN(_01420_));
 OAI21_X1 _26495_ (.A(_16396_),
    .B1(_16344_),
    .B2(_16197_),
    .ZN(_01421_));
 AND3_X1 _26496_ (.A1(_16354_),
    .A2(_16175_),
    .A3(_16367_),
    .ZN(_01422_));
 AOI211_X1 _26497_ (.A(_01422_),
    .B(_16382_),
    .C1(_16302_),
    .C2(_16381_),
    .ZN(_01423_));
 OAI21_X1 _26498_ (.A(_16375_),
    .B1(_16308_),
    .B2(_16399_),
    .ZN(_01424_));
 OAI21_X1 _26499_ (.A(_16381_),
    .B1(_16244_),
    .B2(_16207_),
    .ZN(_01425_));
 AND4_X1 _26500_ (.A1(_16374_),
    .A2(_01423_),
    .A3(_01424_),
    .A4(_01425_),
    .ZN(_01426_));
 NAND2_X1 _26501_ (.A1(_16360_),
    .A2(_16183_),
    .ZN(_01427_));
 OAI21_X1 _26502_ (.A(_16360_),
    .B1(_16257_),
    .B2(_16331_),
    .ZN(_01428_));
 AND4_X1 _26503_ (.A1(_01427_),
    .A2(_16356_),
    .A3(_16363_),
    .A4(_01428_),
    .ZN(_01429_));
 AND2_X1 _26504_ (.A1(_16434_),
    .A2(_16396_),
    .ZN(_01430_));
 AOI211_X1 _26505_ (.A(_01430_),
    .B(_16589_),
    .C1(_01334_),
    .C2(_16396_),
    .ZN(_01431_));
 AND4_X1 _26506_ (.A1(_01421_),
    .A2(_01426_),
    .A3(_01429_),
    .A4(_01431_),
    .ZN(_01432_));
 AOI211_X1 _26507_ (.A(_16649_),
    .B(_16545_),
    .C1(_16508_),
    .C2(_16194_),
    .ZN(_01433_));
 NOR2_X1 _26508_ (.A1(_16389_),
    .A2(_16335_),
    .ZN(_01434_));
 AND2_X1 _26509_ (.A1(_16295_),
    .A2(_16273_),
    .ZN(_01435_));
 AND2_X1 _26510_ (.A1(_16295_),
    .A2(_16377_),
    .ZN(_01436_));
 OR3_X1 _26511_ (.A1(_01434_),
    .A2(_01435_),
    .A3(_01436_),
    .ZN(_01437_));
 AND2_X1 _26512_ (.A1(_16343_),
    .A2(_16339_),
    .ZN(_01438_));
 OR3_X1 _26513_ (.A1(_01438_),
    .A2(_16498_),
    .A3(_16675_),
    .ZN(_01439_));
 AND3_X1 _26514_ (.A1(_16348_),
    .A2(_16171_),
    .A3(_16230_),
    .ZN(_01440_));
 AND2_X1 _26515_ (.A1(_16348_),
    .A2(_16647_),
    .ZN(_01441_));
 NOR4_X1 _26516_ (.A1(_01437_),
    .A2(_01439_),
    .A3(_01440_),
    .A4(_01441_),
    .ZN(_01442_));
 OAI21_X1 _26517_ (.A(_16508_),
    .B1(_16318_),
    .B2(_16624_),
    .ZN(_01443_));
 NAND2_X1 _26518_ (.A1(_16493_),
    .A2(_16377_),
    .ZN(_01444_));
 OAI21_X1 _26519_ (.A(_16305_),
    .B1(_16430_),
    .B2(_16312_),
    .ZN(_01445_));
 AND4_X1 _26520_ (.A1(_01444_),
    .A2(_01386_),
    .A3(_16533_),
    .A4(_01445_),
    .ZN(_01446_));
 AND4_X1 _26521_ (.A1(_01433_),
    .A2(_01442_),
    .A3(_01443_),
    .A4(_01446_),
    .ZN(_01447_));
 NAND2_X1 _26522_ (.A1(_16250_),
    .A2(_16397_),
    .ZN(_01448_));
 NAND4_X1 _26523_ (.A1(_16268_),
    .A2(_16164_),
    .A3(_16167_),
    .A4(_16270_),
    .ZN(_01449_));
 OAI211_X1 _26524_ (.A(_16249_),
    .B(_16198_),
    .C1(_16275_),
    .C2(_16224_),
    .ZN(_01450_));
 AND4_X1 _26525_ (.A1(_01448_),
    .A2(_16548_),
    .A3(_01449_),
    .A4(_01450_),
    .ZN(_01451_));
 NAND3_X1 _26526_ (.A1(_16299_),
    .A2(_16175_),
    .A3(_16268_),
    .ZN(_01452_));
 AND4_X1 _26527_ (.A1(_16429_),
    .A2(_01451_),
    .A3(_16673_),
    .A4(_01452_),
    .ZN(_01453_));
 NAND2_X1 _26528_ (.A1(_16281_),
    .A2(_16354_),
    .ZN(_01454_));
 OAI211_X1 _26529_ (.A(_16281_),
    .B(_16221_),
    .C1(_16239_),
    .C2(_16276_),
    .ZN(_01455_));
 OAI21_X1 _26530_ (.A(_16281_),
    .B1(_16315_),
    .B2(_16434_),
    .ZN(_01456_));
 OAI21_X1 _26531_ (.A(_16280_),
    .B1(_16317_),
    .B2(_16275_),
    .ZN(_01457_));
 AND4_X1 _26532_ (.A1(_01454_),
    .A2(_01455_),
    .A3(_01456_),
    .A4(_01457_),
    .ZN(_01458_));
 OAI21_X1 _26533_ (.A(_16416_),
    .B1(_16357_),
    .B2(_16290_),
    .ZN(_01459_));
 NAND2_X1 _26534_ (.A1(_16416_),
    .A2(_16244_),
    .ZN(_01460_));
 NAND2_X1 _26535_ (.A1(_16416_),
    .A2(_16278_),
    .ZN(_01461_));
 NAND3_X1 _26536_ (.A1(_16207_),
    .A2(_16268_),
    .A3(_16236_),
    .ZN(_01462_));
 AND4_X1 _26537_ (.A1(_16417_),
    .A2(_01460_),
    .A3(_01461_),
    .A4(_01462_),
    .ZN(_01463_));
 AND4_X1 _26538_ (.A1(_01453_),
    .A2(_01458_),
    .A3(_01459_),
    .A4(_01463_),
    .ZN(_01464_));
 NAND4_X1 _26539_ (.A1(_01420_),
    .A2(_01432_),
    .A3(_01447_),
    .A4(_01464_),
    .ZN(_01465_));
 NOR2_X1 _26540_ (.A1(_01465_),
    .A2(_16406_),
    .ZN(_01466_));
 XOR2_X1 _26541_ (.A(_01024_),
    .B(_01023_),
    .Z(_01467_));
 XNOR2_X1 _26542_ (.A(_01466_),
    .B(_01467_),
    .ZN(_01468_));
 MUX2_X1 _26543_ (.A(_01230_),
    .B(_01468_),
    .S(_16040_),
    .Z(_01079_));
 AND2_X1 _26544_ (.A1(_16301_),
    .A2(_16250_),
    .ZN(_01469_));
 OAI211_X1 _26545_ (.A(_16255_),
    .B(_16550_),
    .C1(_16251_),
    .C2(_16625_),
    .ZN(_01470_));
 AOI211_X1 _26546_ (.A(_01469_),
    .B(_01470_),
    .C1(_16258_),
    .C2(_16447_),
    .ZN(_01471_));
 AND4_X1 _26547_ (.A1(_16182_),
    .A2(_16249_),
    .A3(_16193_),
    .A4(_16236_),
    .ZN(_01472_));
 AND2_X1 _26548_ (.A1(_16286_),
    .A2(_16377_),
    .ZN(_01473_));
 AOI211_X1 _26549_ (.A(_01472_),
    .B(_01473_),
    .C1(_16416_),
    .C2(_16194_),
    .ZN(_01474_));
 AND4_X1 _26550_ (.A1(_16569_),
    .A2(_01474_),
    .A3(_01461_),
    .A4(_01462_),
    .ZN(_01475_));
 NAND3_X1 _26551_ (.A1(_16299_),
    .A2(_16225_),
    .A3(_16268_),
    .ZN(_01476_));
 AND2_X1 _26552_ (.A1(_16671_),
    .A2(_01476_),
    .ZN(_01477_));
 AND4_X1 _26553_ (.A1(_16433_),
    .A2(_01477_),
    .A3(_16435_),
    .A4(_01457_),
    .ZN(_01478_));
 AND4_X1 _26554_ (.A1(_16552_),
    .A2(_01393_),
    .A3(_16431_),
    .A4(_01452_),
    .ZN(_01479_));
 AND4_X1 _26555_ (.A1(_01471_),
    .A2(_01475_),
    .A3(_01478_),
    .A4(_01479_),
    .ZN(_01480_));
 AND2_X1 _26556_ (.A1(_16490_),
    .A2(_16187_),
    .ZN(_01481_));
 AND2_X1 _26557_ (.A1(_16357_),
    .A2(_16390_),
    .ZN(_01482_));
 AND3_X1 _26558_ (.A1(_16390_),
    .A2(_16162_),
    .A3(_16221_),
    .ZN(_01483_));
 OR4_X1 _26559_ (.A1(_01481_),
    .A2(_01356_),
    .A3(_01482_),
    .A4(_01483_),
    .ZN(_01484_));
 AOI21_X1 _26560_ (.A(_16369_),
    .B1(_16477_),
    .B2(_16483_),
    .ZN(_01485_));
 NAND2_X1 _26561_ (.A1(_16360_),
    .A2(_16377_),
    .ZN(_01486_));
 NAND4_X1 _26562_ (.A1(_01485_),
    .A2(_16361_),
    .A3(_16364_),
    .A4(_01486_),
    .ZN(_01487_));
 NAND3_X1 _26563_ (.A1(_16220_),
    .A2(_16216_),
    .A3(_16375_),
    .ZN(_01488_));
 NAND2_X1 _26564_ (.A1(_16318_),
    .A2(_16375_),
    .ZN(_01489_));
 OAI211_X1 _26565_ (.A(_01488_),
    .B(_01489_),
    .C1(_16625_),
    .C2(_16379_),
    .ZN(_01490_));
 NAND4_X1 _26566_ (.A1(_16384_),
    .A2(_16480_),
    .A3(_16655_),
    .A4(_16652_),
    .ZN(_01491_));
 NOR4_X1 _26567_ (.A1(_01484_),
    .A2(_01487_),
    .A3(_01490_),
    .A4(_01491_),
    .ZN(_01492_));
 NAND2_X1 _26568_ (.A1(_16178_),
    .A2(_16275_),
    .ZN(_01493_));
 AND3_X1 _26569_ (.A1(_16443_),
    .A2(_01371_),
    .A3(_01493_),
    .ZN(_01494_));
 OAI211_X1 _26570_ (.A(_01494_),
    .B(_16653_),
    .C1(_16260_),
    .C2(_16185_),
    .ZN(_01495_));
 OAI211_X1 _26571_ (.A(_16457_),
    .B(_16426_),
    .C1(_16193_),
    .C2(_16186_),
    .ZN(_01496_));
 OAI211_X1 _26572_ (.A(_01496_),
    .B(_16462_),
    .C1(_16238_),
    .C2(_16622_),
    .ZN(_01497_));
 OAI21_X1 _26573_ (.A(_16582_),
    .B1(_16204_),
    .B2(_16404_),
    .ZN(_01498_));
 OAI21_X1 _26574_ (.A(_16218_),
    .B1(_16207_),
    .B2(_16278_),
    .ZN(_01499_));
 OAI211_X1 _26575_ (.A(_01499_),
    .B(_16641_),
    .C1(_16601_),
    .C2(_16421_),
    .ZN(_01500_));
 NOR4_X1 _26576_ (.A1(_01495_),
    .A2(_01497_),
    .A3(_01498_),
    .A4(_01500_),
    .ZN(_01501_));
 OAI21_X1 _26577_ (.A(_16493_),
    .B1(_16318_),
    .B2(_16624_),
    .ZN(_01502_));
 NAND4_X1 _26578_ (.A1(_16290_),
    .A2(_16424_),
    .A3(_16327_),
    .A4(_16522_),
    .ZN(_01503_));
 NAND4_X1 _26579_ (.A1(_16424_),
    .A2(_16510_),
    .A3(_16239_),
    .A4(_16327_),
    .ZN(_01504_));
 AND3_X1 _26580_ (.A1(_01502_),
    .A2(_01503_),
    .A3(_01504_),
    .ZN(_01505_));
 NOR4_X1 _26581_ (.A1(_16674_),
    .A2(_16646_),
    .A3(_16528_),
    .A4(_01436_),
    .ZN(_01506_));
 AOI21_X1 _26582_ (.A(_16346_),
    .B1(_16419_),
    .B2(_01373_),
    .ZN(_01507_));
 AND3_X1 _26583_ (.A1(_16348_),
    .A2(_16190_),
    .A3(_16164_),
    .ZN(_01508_));
 NOR4_X1 _26584_ (.A1(_01507_),
    .A2(_16497_),
    .A3(_16675_),
    .A4(_01508_),
    .ZN(_01509_));
 AND2_X1 _26585_ (.A1(_16310_),
    .A2(_16322_),
    .ZN(_01510_));
 INV_X1 _26586_ (.A(_01510_),
    .ZN(_01511_));
 NAND3_X1 _26587_ (.A1(_16508_),
    .A2(_16171_),
    .A3(_16230_),
    .ZN(_01512_));
 OAI21_X1 _26588_ (.A(_16508_),
    .B1(_16357_),
    .B2(_16344_),
    .ZN(_01513_));
 AND4_X1 _26589_ (.A1(_16323_),
    .A2(_01511_),
    .A3(_01512_),
    .A4(_01513_),
    .ZN(_01514_));
 AND4_X1 _26590_ (.A1(_01505_),
    .A2(_01506_),
    .A3(_01509_),
    .A4(_01514_),
    .ZN(_01515_));
 NAND4_X1 _26591_ (.A1(_01480_),
    .A2(_01492_),
    .A3(_01501_),
    .A4(_01515_),
    .ZN(_01516_));
 NOR2_X1 _26592_ (.A1(_01516_),
    .A2(_16406_),
    .ZN(_01517_));
 XOR2_X1 _26593_ (.A(_01026_),
    .B(_01025_),
    .Z(_01518_));
 XNOR2_X1 _26594_ (.A(_01517_),
    .B(_01518_),
    .ZN(_01519_));
 MUX2_X1 _26595_ (.A(_01231_),
    .B(_01519_),
    .S(_16040_),
    .Z(_01081_));
 AND2_X1 _26596_ (.A1(_16258_),
    .A2(_16306_),
    .ZN(_01520_));
 AOI211_X1 _26597_ (.A(_01520_),
    .B(_01469_),
    .C1(_16430_),
    .C2(_16258_),
    .ZN(_01521_));
 OAI211_X1 _26598_ (.A(_16424_),
    .B(_16269_),
    .C1(_16197_),
    .C2(_16486_),
    .ZN(_01522_));
 OAI211_X1 _26599_ (.A(_16424_),
    .B(_16269_),
    .C1(_16275_),
    .C2(_16483_),
    .ZN(_01523_));
 AND4_X1 _26600_ (.A1(_16673_),
    .A2(_01521_),
    .A3(_01522_),
    .A4(_01523_),
    .ZN(_01524_));
 AND2_X1 _26601_ (.A1(_16283_),
    .A2(_16348_),
    .ZN(_01525_));
 AND2_X1 _26602_ (.A1(_16265_),
    .A2(_16348_),
    .ZN(_01526_));
 OR4_X1 _26603_ (.A1(_16498_),
    .A2(_01525_),
    .A3(_01526_),
    .A4(_01441_),
    .ZN(_01527_));
 OAI21_X1 _26604_ (.A(_16643_),
    .B1(_16335_),
    .B2(_16378_),
    .ZN(_01528_));
 AOI21_X1 _26605_ (.A(_16335_),
    .B1(_01336_),
    .B2(_16421_),
    .ZN(_01529_));
 OAI21_X1 _26606_ (.A(_16502_),
    .B1(_16168_),
    .B2(_16335_),
    .ZN(_01530_));
 NOR4_X1 _26607_ (.A1(_01527_),
    .A2(_01528_),
    .A3(_01529_),
    .A4(_01530_),
    .ZN(_01531_));
 NAND3_X1 _26608_ (.A1(_16308_),
    .A2(_16424_),
    .A3(_16327_),
    .ZN(_01532_));
 OAI211_X1 _26609_ (.A(_16424_),
    .B(_16327_),
    .C1(_16275_),
    .C2(_16278_),
    .ZN(_01533_));
 NAND4_X1 _26610_ (.A1(_16664_),
    .A2(_01386_),
    .A3(_01532_),
    .A4(_01533_),
    .ZN(_01534_));
 AOI211_X1 _26611_ (.A(_16234_),
    .B(_16540_),
    .C1(_16239_),
    .C2(_16276_),
    .ZN(_01535_));
 AOI21_X1 _26612_ (.A(_16540_),
    .B1(_16300_),
    .B2(_16191_),
    .ZN(_01536_));
 NOR4_X1 _26613_ (.A1(_01534_),
    .A2(_01510_),
    .A3(_01535_),
    .A4(_01536_),
    .ZN(_01537_));
 OAI21_X1 _26614_ (.A(_16281_),
    .B1(_16317_),
    .B2(_16278_),
    .ZN(_01538_));
 NAND4_X1 _26615_ (.A1(_01538_),
    .A2(_16433_),
    .A3(_16566_),
    .A4(_01476_),
    .ZN(_01539_));
 NAND2_X1 _26616_ (.A1(_16417_),
    .A2(_01462_),
    .ZN(_01540_));
 NOR4_X1 _26617_ (.A1(_01539_),
    .A2(_01540_),
    .A3(_16287_),
    .A4(_01473_),
    .ZN(_01541_));
 NAND4_X1 _26618_ (.A1(_01524_),
    .A2(_01531_),
    .A3(_01537_),
    .A4(_01541_),
    .ZN(_01542_));
 AND2_X1 _26619_ (.A1(_16385_),
    .A2(_16306_),
    .ZN(_01543_));
 AOI211_X1 _26620_ (.A(_01422_),
    .B(_01543_),
    .C1(_16385_),
    .C2(_16486_),
    .ZN(_01544_));
 OAI21_X1 _26621_ (.A(_16385_),
    .B1(_16414_),
    .B2(_16275_),
    .ZN(_01545_));
 OAI21_X1 _26622_ (.A(_16375_),
    .B1(_16357_),
    .B2(_16344_),
    .ZN(_01546_));
 OAI21_X1 _26623_ (.A(_16375_),
    .B1(_16207_),
    .B2(_16331_),
    .ZN(_01547_));
 AND4_X1 _26624_ (.A1(_01544_),
    .A2(_01545_),
    .A3(_01546_),
    .A4(_01547_),
    .ZN(_01548_));
 NAND2_X1 _26625_ (.A1(_01412_),
    .A2(_16180_),
    .ZN(_01549_));
 OAI211_X1 _26626_ (.A(_01549_),
    .B(_16446_),
    .C1(_16544_),
    .C2(_16185_),
    .ZN(_01550_));
 NAND4_X1 _26627_ (.A1(_16445_),
    .A2(_16577_),
    .A3(_16575_),
    .A4(_01493_),
    .ZN(_01551_));
 AND3_X1 _26628_ (.A1(_16617_),
    .A2(_16522_),
    .A3(_16450_),
    .ZN(_01552_));
 AOI211_X1 _26629_ (.A(_16234_),
    .B(_16204_),
    .C1(_10987_),
    .C2(_10993_),
    .ZN(_01553_));
 NOR4_X1 _26630_ (.A1(_01550_),
    .A2(_01551_),
    .A3(_01552_),
    .A4(_01553_),
    .ZN(_01554_));
 OAI21_X1 _26631_ (.A(_16477_),
    .B1(_16283_),
    .B2(_16228_),
    .ZN(_01555_));
 NAND4_X1 _26632_ (.A1(_16359_),
    .A2(_01427_),
    .A3(_01486_),
    .A4(_01555_),
    .ZN(_01556_));
 NAND2_X1 _26633_ (.A1(_16302_),
    .A2(_16396_),
    .ZN(_01557_));
 NAND2_X1 _26634_ (.A1(_16357_),
    .A2(_16396_),
    .ZN(_01558_));
 NAND3_X1 _26635_ (.A1(_01557_),
    .A2(_01558_),
    .A3(_16487_),
    .ZN(_01559_));
 NOR4_X1 _26636_ (.A1(_01556_),
    .A2(_01357_),
    .A3(_01481_),
    .A4(_01559_),
    .ZN(_01560_));
 OAI21_X1 _26637_ (.A(_16457_),
    .B1(_16207_),
    .B2(_16647_),
    .ZN(_01561_));
 OAI21_X1 _26638_ (.A(_16219_),
    .B1(_16232_),
    .B2(_16318_),
    .ZN(_01562_));
 OAI21_X1 _26639_ (.A(_16219_),
    .B1(_16197_),
    .B2(_16265_),
    .ZN(_01563_));
 OAI211_X1 _26640_ (.A(_16457_),
    .B(_10987_),
    .C1(_16510_),
    .C2(_16221_),
    .ZN(_01564_));
 AND4_X1 _26641_ (.A1(_01561_),
    .A2(_01562_),
    .A3(_01563_),
    .A4(_01564_),
    .ZN(_01565_));
 NAND4_X1 _26642_ (.A1(_01548_),
    .A2(_01554_),
    .A3(_01560_),
    .A4(_01565_),
    .ZN(_01566_));
 NOR2_X1 _26643_ (.A1(_01542_),
    .A2(_01566_),
    .ZN(_01567_));
 XOR2_X1 _26644_ (.A(_01028_),
    .B(_01027_),
    .Z(_01568_));
 XNOR2_X1 _26645_ (.A(_01567_),
    .B(_01568_),
    .ZN(_01569_));
 BUF_X2 _26646_ (.A(_03738_),
    .Z(_01570_));
 MUX2_X1 _26647_ (.A(_01232_),
    .B(_01569_),
    .S(_01570_),
    .Z(_01082_));
 XOR2_X1 _26648_ (.A(_17165_),
    .B(_17000_),
    .Z(_01571_));
 XNOR2_X1 _26649_ (.A(_13842_),
    .B(_12727_),
    .ZN(_01572_));
 XNOR2_X1 _26650_ (.A(_01572_),
    .B(_13287_),
    .ZN(_01573_));
 XNOR2_X1 _26651_ (.A(_13019_),
    .B(_01573_),
    .ZN(_01574_));
 XNOR2_X1 _26652_ (.A(_01574_),
    .B(_17165_),
    .ZN(_01575_));
 MUX2_X1 _26653_ (.A(_01571_),
    .B(_01575_),
    .S(_15155_),
    .Z(_00687_));
 XOR2_X1 _26654_ (.A(_17166_),
    .B(_17001_),
    .Z(_01576_));
 XOR2_X1 _26655_ (.A(_13288_),
    .B(_13515_),
    .Z(_01577_));
 XOR2_X2 _26656_ (.A(_13842_),
    .B(_13094_),
    .Z(_01578_));
 XNOR2_X1 _26657_ (.A(_13217_),
    .B(_01578_),
    .ZN(_01579_));
 XNOR2_X1 _26658_ (.A(_01577_),
    .B(_01579_),
    .ZN(_01580_));
 XNOR2_X1 _26659_ (.A(_01580_),
    .B(_17166_),
    .ZN(_01581_));
 MUX2_X1 _26660_ (.A(_01576_),
    .B(_01581_),
    .S(_15155_),
    .Z(_00688_));
 XOR2_X1 _26661_ (.A(_17167_),
    .B(_17002_),
    .Z(_01582_));
 XNOR2_X1 _26662_ (.A(_13791_),
    .B(_13346_),
    .ZN(_01583_));
 XNOR2_X1 _26663_ (.A(_13516_),
    .B(_01583_),
    .ZN(_01584_));
 XOR2_X1 _26664_ (.A(_01584_),
    .B(_17167_),
    .Z(_01585_));
 MUX2_X1 _26665_ (.A(_01582_),
    .B(_01585_),
    .S(_15155_),
    .Z(_00689_));
 XOR2_X1 _26666_ (.A(_17168_),
    .B(_17003_),
    .Z(_01586_));
 XOR2_X2 _26667_ (.A(_13791_),
    .B(_13580_),
    .Z(_01587_));
 XNOR2_X1 _26668_ (.A(_01587_),
    .B(_13686_),
    .ZN(_01588_));
 XNOR2_X1 _26669_ (.A(_01588_),
    .B(_13946_),
    .ZN(_01589_));
 XOR2_X1 _26670_ (.A(_01589_),
    .B(_17168_),
    .Z(_01590_));
 MUX2_X1 _26671_ (.A(_01586_),
    .B(_01590_),
    .S(_15155_),
    .Z(_00690_));
 XOR2_X1 _26672_ (.A(_17169_),
    .B(_17004_),
    .Z(_01591_));
 XNOR2_X1 _26673_ (.A(_13946_),
    .B(_13736_),
    .ZN(_01592_));
 XNOR2_X1 _26674_ (.A(_01592_),
    .B(_13896_),
    .ZN(_01593_));
 XNOR2_X1 _26675_ (.A(_01593_),
    .B(_12101_),
    .ZN(_01594_));
 XNOR2_X1 _26676_ (.A(_01594_),
    .B(_17169_),
    .ZN(_01595_));
 MUX2_X1 _26677_ (.A(_01591_),
    .B(_01595_),
    .S(_15155_),
    .Z(_00691_));
 XOR2_X2 _26678_ (.A(_17131_),
    .B(_17099_),
    .Z(_01596_));
 XNOR2_X1 _26679_ (.A(_14165_),
    .B(_01596_),
    .ZN(_01597_));
 MUX2_X1 _26680_ (.A(_01290_),
    .B(_01597_),
    .S(_01570_),
    .Z(_01090_));
 XOR2_X1 _26681_ (.A(_17142_),
    .B(_17110_),
    .Z(_01598_));
 XNOR2_X1 _26682_ (.A(_14283_),
    .B(_01598_),
    .ZN(_01599_));
 MUX2_X1 _26683_ (.A(_01291_),
    .B(_01599_),
    .S(_01570_),
    .Z(_01101_));
 XOR2_X2 _26684_ (.A(_17153_),
    .B(_17121_),
    .Z(_01600_));
 XNOR2_X1 _26685_ (.A(_14368_),
    .B(_01600_),
    .ZN(_01601_));
 MUX2_X1 _26686_ (.A(_01292_),
    .B(_01601_),
    .S(_01570_),
    .Z(_01112_));
 XOR2_X2 _26687_ (.A(_17156_),
    .B(_17124_),
    .Z(_01602_));
 XNOR2_X2 _26688_ (.A(_14439_),
    .B(_01602_),
    .ZN(_01603_));
 MUX2_X1 _26689_ (.A(_01293_),
    .B(_01603_),
    .S(_01570_),
    .Z(_01115_));
 AND2_X1 _26690_ (.A1(_14467_),
    .A2(_14490_),
    .ZN(_01604_));
 XOR2_X2 _26691_ (.A(_17157_),
    .B(_17125_),
    .Z(_01605_));
 XNOR2_X1 _26692_ (.A(_01604_),
    .B(_01605_),
    .ZN(_01606_));
 MUX2_X1 _26693_ (.A(_01294_),
    .B(_01606_),
    .S(_01570_),
    .Z(_01116_));
 XOR2_X2 _26694_ (.A(_17158_),
    .B(_17126_),
    .Z(_01607_));
 XNOR2_X1 _26695_ (.A(_14554_),
    .B(_01607_),
    .ZN(_01608_));
 MUX2_X1 _26696_ (.A(_01295_),
    .B(_01608_),
    .S(_01570_),
    .Z(_01117_));
 XOR2_X1 _26697_ (.A(_17159_),
    .B(_17127_),
    .Z(_01609_));
 XNOR2_X1 _26698_ (.A(_14610_),
    .B(_01609_),
    .ZN(_01610_));
 MUX2_X1 _26699_ (.A(_01297_),
    .B(_01610_),
    .S(_01570_),
    .Z(_01118_));
 XOR2_X2 _26700_ (.A(_17160_),
    .B(_17128_),
    .Z(_01611_));
 XNOR2_X1 _26701_ (.A(_14659_),
    .B(_01611_),
    .ZN(_01612_));
 MUX2_X1 _26702_ (.A(_01298_),
    .B(_01612_),
    .S(_01570_),
    .Z(_01119_));
 XOR2_X2 _26703_ (.A(_17161_),
    .B(_17129_),
    .Z(_01613_));
 XNOR2_X1 _26704_ (.A(_14876_),
    .B(_01613_),
    .ZN(_01614_));
 MUX2_X1 _26705_ (.A(_01299_),
    .B(_01614_),
    .S(_01570_),
    .Z(_01120_));
 NOR2_X1 _26706_ (.A1(_03749_),
    .A2(_01300_),
    .ZN(_01615_));
 XNOR2_X1 _26707_ (.A(_17162_),
    .B(_17130_),
    .ZN(_01616_));
 XNOR2_X1 _26708_ (.A(_14976_),
    .B(_01616_),
    .ZN(_01617_));
 AOI21_X1 _26709_ (.A(_01615_),
    .B1(_01617_),
    .B2(_03749_),
    .ZN(_01121_));
 XOR2_X2 _26710_ (.A(_17132_),
    .B(_17100_),
    .Z(_01618_));
 XNOR2_X1 _26711_ (.A(_15064_),
    .B(_01618_),
    .ZN(_01619_));
 BUF_X2 _26712_ (.A(_03738_),
    .Z(_01620_));
 MUX2_X1 _26713_ (.A(_01301_),
    .B(_01619_),
    .S(_01620_),
    .Z(_01091_));
 XOR2_X2 _26714_ (.A(_17133_),
    .B(_17101_),
    .Z(_01621_));
 XNOR2_X1 _26715_ (.A(_15145_),
    .B(_01621_),
    .ZN(_01622_));
 MUX2_X1 _26716_ (.A(_01302_),
    .B(_01622_),
    .S(_01620_),
    .Z(_01092_));
 XOR2_X2 _26717_ (.A(_17134_),
    .B(_17102_),
    .Z(_01623_));
 XNOR2_X1 _26718_ (.A(_15212_),
    .B(_01623_),
    .ZN(_01624_));
 MUX2_X1 _26719_ (.A(_01303_),
    .B(_01624_),
    .S(_01620_),
    .Z(_01093_));
 XOR2_X2 _26720_ (.A(_17135_),
    .B(_17103_),
    .Z(_01625_));
 XNOR2_X1 _26721_ (.A(_15283_),
    .B(_01625_),
    .ZN(_01626_));
 MUX2_X1 _26722_ (.A(_01304_),
    .B(_01626_),
    .S(_01620_),
    .Z(_01094_));
 XOR2_X2 _26723_ (.A(_17136_),
    .B(_17104_),
    .Z(_01627_));
 XNOR2_X1 _26724_ (.A(_15345_),
    .B(_01627_),
    .ZN(_01628_));
 MUX2_X1 _26725_ (.A(_01305_),
    .B(_01628_),
    .S(_01620_),
    .Z(_01095_));
 XOR2_X2 _26726_ (.A(_17137_),
    .B(_17105_),
    .Z(_01629_));
 XNOR2_X1 _26727_ (.A(_15405_),
    .B(_01629_),
    .ZN(_01630_));
 MUX2_X1 _26728_ (.A(_01306_),
    .B(_01630_),
    .S(_01620_),
    .Z(_01096_));
 XOR2_X1 _26729_ (.A(_17138_),
    .B(_17106_),
    .Z(_01631_));
 XNOR2_X1 _26730_ (.A(_15642_),
    .B(_01631_),
    .ZN(_01632_));
 MUX2_X1 _26731_ (.A(_01308_),
    .B(_01632_),
    .S(_01620_),
    .Z(_01097_));
 NAND2_X1 _26732_ (.A1(_03847_),
    .A2(_01309_),
    .ZN(_01633_));
 XOR2_X1 _26733_ (.A(_17139_),
    .B(_17107_),
    .Z(_01634_));
 XOR2_X1 _26734_ (.A(_15748_),
    .B(_01634_),
    .Z(_01635_));
 OAI21_X1 _26735_ (.A(_01633_),
    .B1(_01635_),
    .B2(_03847_),
    .ZN(_01098_));
 XOR2_X1 _26736_ (.A(_17140_),
    .B(_17108_),
    .Z(_01636_));
 XNOR2_X1 _26737_ (.A(_15832_),
    .B(_01636_),
    .ZN(_01637_));
 MUX2_X1 _26738_ (.A(_01310_),
    .B(_01637_),
    .S(_01620_),
    .Z(_01099_));
 XOR2_X1 _26739_ (.A(_17141_),
    .B(_17109_),
    .Z(_01638_));
 XNOR2_X1 _26740_ (.A(_15911_),
    .B(_01638_),
    .ZN(_01639_));
 MUX2_X1 _26741_ (.A(_01311_),
    .B(_01639_),
    .S(_01620_),
    .Z(_01100_));
 XOR2_X1 _26742_ (.A(_17143_),
    .B(_17111_),
    .Z(_01640_));
 XNOR2_X1 _26743_ (.A(_15974_),
    .B(_01640_),
    .ZN(_01641_));
 MUX2_X1 _26744_ (.A(_01312_),
    .B(_01641_),
    .S(_01620_),
    .Z(_01102_));
 NOR2_X1 _26745_ (.A1(_03749_),
    .A2(_01313_),
    .ZN(_01642_));
 XOR2_X1 _26746_ (.A(_17144_),
    .B(_17112_),
    .Z(_01643_));
 XOR2_X1 _26747_ (.A(_16038_),
    .B(_01643_),
    .Z(_01644_));
 AOI21_X1 _26748_ (.A(_01642_),
    .B1(_01644_),
    .B2(_03749_),
    .ZN(_01103_));
 NAND2_X1 _26749_ (.A1(_03847_),
    .A2(_01314_),
    .ZN(_01645_));
 XOR2_X1 _26750_ (.A(_17145_),
    .B(_17113_),
    .Z(_01646_));
 XOR2_X1 _26751_ (.A(_16110_),
    .B(_01646_),
    .Z(_01647_));
 OAI21_X1 _26752_ (.A(_01645_),
    .B1(_01647_),
    .B2(_03847_),
    .ZN(_01104_));
 XOR2_X1 _26753_ (.A(_17146_),
    .B(_17114_),
    .Z(_01648_));
 XNOR2_X1 _26754_ (.A(_16160_),
    .B(_01648_),
    .ZN(_01649_));
 BUF_X2 _26755_ (.A(_03933_),
    .Z(_01650_));
 MUX2_X1 _26756_ (.A(_01315_),
    .B(_01649_),
    .S(_01650_),
    .Z(_01105_));
 XNOR2_X1 _26757_ (.A(_01013_),
    .B(_17115_),
    .ZN(_01651_));
 XNOR2_X1 _26758_ (.A(_01651_),
    .B(_17147_),
    .ZN(_01652_));
 XNOR2_X1 _26759_ (.A(_16408_),
    .B(_01652_),
    .ZN(_01653_));
 MUX2_X1 _26760_ (.A(_01316_),
    .B(_01653_),
    .S(_01650_),
    .Z(_01106_));
 XOR2_X1 _26761_ (.A(_01015_),
    .B(_17116_),
    .Z(_01654_));
 XNOR2_X1 _26762_ (.A(_01654_),
    .B(_17148_),
    .ZN(_01655_));
 XNOR2_X1 _26763_ (.A(_16518_),
    .B(_01655_),
    .ZN(_01656_));
 MUX2_X1 _26764_ (.A(_01317_),
    .B(_01656_),
    .S(_01650_),
    .Z(_01107_));
 XNOR2_X1 _26765_ (.A(_01017_),
    .B(_17117_),
    .ZN(_01657_));
 INV_X1 _26766_ (.A(_17149_),
    .ZN(_01658_));
 XNOR2_X1 _26767_ (.A(_01657_),
    .B(_01658_),
    .ZN(_01659_));
 XNOR2_X1 _26768_ (.A(_16608_),
    .B(_01659_),
    .ZN(_01660_));
 MUX2_X1 _26769_ (.A(_01319_),
    .B(_01660_),
    .S(_01650_),
    .Z(_01108_));
 XNOR2_X1 _26770_ (.A(_01019_),
    .B(_17118_),
    .ZN(_01661_));
 INV_X1 _26771_ (.A(_17150_),
    .ZN(_01662_));
 XNOR2_X1 _26772_ (.A(_01661_),
    .B(_01662_),
    .ZN(_01663_));
 XNOR2_X1 _26773_ (.A(_01341_),
    .B(_01663_),
    .ZN(_01664_));
 MUX2_X1 _26774_ (.A(_01320_),
    .B(_01664_),
    .S(_01650_),
    .Z(_01109_));
 XOR2_X1 _26775_ (.A(_01021_),
    .B(_17119_),
    .Z(_01665_));
 XNOR2_X1 _26776_ (.A(_01665_),
    .B(_17151_),
    .ZN(_01666_));
 XNOR2_X1 _26777_ (.A(_01404_),
    .B(_01666_),
    .ZN(_01667_));
 MUX2_X1 _26778_ (.A(_01321_),
    .B(_01667_),
    .S(_01650_),
    .Z(_01110_));
 XOR2_X1 _26779_ (.A(_01023_),
    .B(_17120_),
    .Z(_01668_));
 XNOR2_X1 _26780_ (.A(_01668_),
    .B(_17152_),
    .ZN(_01669_));
 XNOR2_X1 _26781_ (.A(_01466_),
    .B(_01669_),
    .ZN(_01670_));
 MUX2_X1 _26782_ (.A(_01322_),
    .B(_01670_),
    .S(_01650_),
    .Z(_01111_));
 XOR2_X1 _26783_ (.A(_01025_),
    .B(_17122_),
    .Z(_01671_));
 XNOR2_X1 _26784_ (.A(_01671_),
    .B(_17154_),
    .ZN(_01672_));
 XNOR2_X1 _26785_ (.A(_01517_),
    .B(_01672_),
    .ZN(_01673_));
 MUX2_X1 _26786_ (.A(_01323_),
    .B(_01673_),
    .S(_01650_),
    .Z(_01113_));
 XOR2_X1 _26787_ (.A(_01027_),
    .B(_17123_),
    .Z(_01674_));
 XNOR2_X1 _26788_ (.A(_01674_),
    .B(_17155_),
    .ZN(_01675_));
 XNOR2_X1 _26789_ (.A(_01567_),
    .B(_01675_),
    .ZN(_01676_));
 MUX2_X1 _26790_ (.A(_01324_),
    .B(_01676_),
    .S(_01650_),
    .Z(_01114_));
 XOR2_X1 _26791_ (.A(_17170_),
    .B(_17005_),
    .Z(_01677_));
 XNOR2_X1 _26792_ (.A(_13895_),
    .B(_01029_),
    .ZN(_01678_));
 XOR2_X1 _26793_ (.A(_15149_),
    .B(_01678_),
    .Z(_01679_));
 XOR2_X1 _26794_ (.A(_12499_),
    .B(_11776_),
    .Z(_01680_));
 XNOR2_X1 _26795_ (.A(_01679_),
    .B(_01680_),
    .ZN(_01681_));
 MUX2_X1 _26796_ (.A(_01677_),
    .B(_01681_),
    .S(_15155_),
    .Z(_00652_));
 XOR2_X1 _26797_ (.A(_17171_),
    .B(_17006_),
    .Z(_01682_));
 XNOR2_X1 _26798_ (.A(_12181_),
    .B(_01030_),
    .ZN(_01683_));
 XNOR2_X1 _26799_ (.A(_11312_),
    .B(_13895_),
    .ZN(_01684_));
 XNOR2_X1 _26800_ (.A(_01683_),
    .B(_01684_),
    .ZN(_01685_));
 XNOR2_X1 _26801_ (.A(_16042_),
    .B(_15149_),
    .ZN(_01686_));
 XNOR2_X1 _26802_ (.A(_01685_),
    .B(_01686_),
    .ZN(_01687_));
 MUX2_X1 _26803_ (.A(_01682_),
    .B(_01687_),
    .S(_15155_),
    .Z(_00653_));
 XOR2_X1 _26804_ (.A(_12727_),
    .B(_12575_),
    .Z(_01688_));
 XNOR2_X1 _26805_ (.A(_01688_),
    .B(_13017_),
    .ZN(_01689_));
 XNOR2_X1 _26806_ (.A(_12385_),
    .B(_12284_),
    .ZN(_01690_));
 OAI21_X1 _26807_ (.A(_09038_),
    .B1(_01689_),
    .B2(_01690_),
    .ZN(_01691_));
 AOI21_X1 _26808_ (.A(_01691_),
    .B1(_01689_),
    .B2(_01690_),
    .ZN(_01692_));
 AND2_X1 _26809_ (.A1(_01331_),
    .A2(_17008_),
    .ZN(_01693_));
 NOR2_X1 _26810_ (.A1(_01692_),
    .A2(_01693_),
    .ZN(_01694_));
 XNOR2_X1 _26811_ (.A(_01694_),
    .B(_17172_),
    .ZN(_00654_));
 XOR2_X1 _26812_ (.A(_17173_),
    .B(_17009_),
    .Z(_01695_));
 XNOR2_X1 _26813_ (.A(_13287_),
    .B(_12727_),
    .ZN(_01696_));
 XNOR2_X1 _26814_ (.A(_01696_),
    .B(_01578_),
    .ZN(_01697_));
 XOR2_X2 _26815_ (.A(_13895_),
    .B(_12650_),
    .Z(_01698_));
 XNOR2_X1 _26816_ (.A(_01698_),
    .B(_12952_),
    .ZN(_01699_));
 XNOR2_X1 _26817_ (.A(_01697_),
    .B(_01699_),
    .ZN(_01700_));
 XNOR2_X1 _26818_ (.A(_01700_),
    .B(_17173_),
    .ZN(_01701_));
 MUX2_X1 _26819_ (.A(_01695_),
    .B(_01701_),
    .S(_15155_),
    .Z(_00655_));
 XOR2_X1 _26820_ (.A(_17175_),
    .B(_17010_),
    .Z(_01702_));
 XNOR2_X1 _26821_ (.A(_12883_),
    .B(_13895_),
    .ZN(_01703_));
 XOR2_X1 _26822_ (.A(_01703_),
    .B(_13159_),
    .Z(_01704_));
 XNOR2_X1 _26823_ (.A(_01578_),
    .B(_13346_),
    .ZN(_01705_));
 XNOR2_X1 _26824_ (.A(_01704_),
    .B(_01705_),
    .ZN(_01706_));
 XNOR2_X1 _26825_ (.A(_01706_),
    .B(_13515_),
    .ZN(_01707_));
 INV_X1 _26826_ (.A(_17175_),
    .ZN(_01708_));
 XNOR2_X1 _26827_ (.A(_01707_),
    .B(_01708_),
    .ZN(_01709_));
 BUF_X2 _26828_ (.A(_09039_),
    .Z(_01710_));
 MUX2_X1 _26829_ (.A(_01702_),
    .B(_01709_),
    .S(_01710_),
    .Z(_00656_));
 XOR2_X1 _26830_ (.A(_17176_),
    .B(_17011_),
    .Z(_01711_));
 XNOR2_X1 _26831_ (.A(_01587_),
    .B(_13216_),
    .ZN(_01712_));
 XNOR2_X1 _26832_ (.A(_13346_),
    .B(_01031_),
    .ZN(_01713_));
 XNOR2_X1 _26833_ (.A(_01713_),
    .B(_13463_),
    .ZN(_01714_));
 XNOR2_X1 _26834_ (.A(_01712_),
    .B(_01714_),
    .ZN(_01715_));
 MUX2_X1 _26835_ (.A(_01711_),
    .B(_01715_),
    .S(_01710_),
    .Z(_00657_));
 XOR2_X1 _26836_ (.A(_17177_),
    .B(_17012_),
    .Z(_01716_));
 XNOR2_X1 _26837_ (.A(_13736_),
    .B(_01032_),
    .ZN(_01717_));
 XOR2_X1 _26838_ (.A(_01717_),
    .B(_13408_),
    .Z(_01718_));
 XNOR2_X1 _26839_ (.A(_13685_),
    .B(_13580_),
    .ZN(_01719_));
 XNOR2_X1 _26840_ (.A(_01719_),
    .B(_13946_),
    .ZN(_01720_));
 XNOR2_X1 _26841_ (.A(_01718_),
    .B(_01720_),
    .ZN(_01721_));
 MUX2_X1 _26842_ (.A(_01716_),
    .B(_01721_),
    .S(_01710_),
    .Z(_00658_));
 XOR2_X1 _26843_ (.A(_17178_),
    .B(_17013_),
    .Z(_01722_));
 XOR2_X1 _26844_ (.A(_13736_),
    .B(_11877_),
    .Z(_01723_));
 XNOR2_X1 _26845_ (.A(_13637_),
    .B(_13842_),
    .ZN(_01724_));
 XNOR2_X1 _26846_ (.A(_01723_),
    .B(_01724_),
    .ZN(_01725_));
 XNOR2_X1 _26847_ (.A(_01725_),
    .B(_12101_),
    .ZN(_01726_));
 INV_X1 _26848_ (.A(_17178_),
    .ZN(_01727_));
 XNOR2_X1 _26849_ (.A(_01726_),
    .B(_01727_),
    .ZN(_01728_));
 MUX2_X1 _26850_ (.A(_01722_),
    .B(_01728_),
    .S(_01710_),
    .Z(_00659_));
 XOR2_X1 _26851_ (.A(_01597_),
    .B(_17163_),
    .Z(_01729_));
 MUX2_X1 _26852_ (.A(_01255_),
    .B(_01729_),
    .S(_01650_),
    .Z(_01122_));
 INV_X1 _26853_ (.A(_17174_),
    .ZN(_01730_));
 MUX2_X1 _26854_ (.A(_17174_),
    .B(_01256_),
    .S(_01330_),
    .Z(_01731_));
 NAND2_X1 _26855_ (.A1(_01599_),
    .A2(_03738_),
    .ZN(_01732_));
 MUX2_X1 _26856_ (.A(_01730_),
    .B(_01731_),
    .S(_01732_),
    .Z(_01133_));
 INV_X1 _26857_ (.A(_17185_),
    .ZN(_01733_));
 XNOR2_X1 _26858_ (.A(_01601_),
    .B(_01733_),
    .ZN(_01734_));
 BUF_X2 _26859_ (.A(_03933_),
    .Z(_01735_));
 MUX2_X1 _26860_ (.A(_01257_),
    .B(_01734_),
    .S(_01735_),
    .Z(_01144_));
 BUF_X2 _26861_ (.A(_03933_),
    .Z(_01736_));
 AND3_X1 _26862_ (.A1(_01603_),
    .A2(_01736_),
    .A3(_17188_),
    .ZN(_01737_));
 MUX2_X1 _26863_ (.A(_17188_),
    .B(_01258_),
    .S(_01330_),
    .Z(_01738_));
 AOI21_X1 _26864_ (.A(_01738_),
    .B1(_01603_),
    .B2(_03749_),
    .ZN(_01739_));
 NOR2_X1 _26865_ (.A1(_01737_),
    .A2(_01739_),
    .ZN(_01147_));
 XNOR2_X1 _26866_ (.A(_01605_),
    .B(_17189_),
    .ZN(_01740_));
 XOR2_X1 _26867_ (.A(_01604_),
    .B(_01740_),
    .Z(_01741_));
 MUX2_X1 _26868_ (.A(_01259_),
    .B(_01741_),
    .S(_01735_),
    .Z(_01148_));
 INV_X1 _26869_ (.A(_17190_),
    .ZN(_01742_));
 XNOR2_X1 _26870_ (.A(_01608_),
    .B(_01742_),
    .ZN(_01743_));
 MUX2_X1 _26871_ (.A(_01260_),
    .B(_01743_),
    .S(_01735_),
    .Z(_01149_));
 XOR2_X1 _26872_ (.A(_17191_),
    .B(_17159_),
    .Z(_01744_));
 XOR2_X1 _26873_ (.A(_01744_),
    .B(_17127_),
    .Z(_01745_));
 XNOR2_X1 _26874_ (.A(_14610_),
    .B(_01745_),
    .ZN(_01746_));
 MUX2_X1 _26875_ (.A(_01261_),
    .B(_01746_),
    .S(_01735_),
    .Z(_01150_));
 XNOR2_X1 _26876_ (.A(_01611_),
    .B(_17192_),
    .ZN(_01747_));
 XOR2_X1 _26877_ (.A(_14659_),
    .B(_01747_),
    .Z(_01748_));
 MUX2_X1 _26878_ (.A(_01262_),
    .B(_01748_),
    .S(_01735_),
    .Z(_01151_));
 XNOR2_X1 _26879_ (.A(_01613_),
    .B(_17193_),
    .ZN(_01749_));
 XOR2_X1 _26880_ (.A(_14876_),
    .B(_01749_),
    .Z(_01750_));
 MUX2_X1 _26881_ (.A(_01264_),
    .B(_01750_),
    .S(_01735_),
    .Z(_01152_));
 XNOR2_X1 _26882_ (.A(_01616_),
    .B(_15153_),
    .ZN(_01751_));
 XOR2_X1 _26883_ (.A(_14976_),
    .B(_01751_),
    .Z(_01752_));
 MUX2_X1 _26884_ (.A(_01265_),
    .B(_01752_),
    .S(_01735_),
    .Z(_01153_));
 XOR2_X1 _26885_ (.A(_01619_),
    .B(_17164_),
    .Z(_01753_));
 MUX2_X1 _26886_ (.A(_01266_),
    .B(_01753_),
    .S(_01735_),
    .Z(_01123_));
 XOR2_X1 _26887_ (.A(_01622_),
    .B(_17165_),
    .Z(_01754_));
 MUX2_X1 _26888_ (.A(_01267_),
    .B(_01754_),
    .S(_01735_),
    .Z(_01124_));
 INV_X1 _26889_ (.A(_17166_),
    .ZN(_01755_));
 XNOR2_X1 _26890_ (.A(_01624_),
    .B(_01755_),
    .ZN(_01756_));
 MUX2_X1 _26891_ (.A(_01268_),
    .B(_01756_),
    .S(_01735_),
    .Z(_01125_));
 XOR2_X1 _26892_ (.A(_01626_),
    .B(_17167_),
    .Z(_01757_));
 BUF_X2 _26893_ (.A(_03933_),
    .Z(_01758_));
 MUX2_X1 _26894_ (.A(_01269_),
    .B(_01757_),
    .S(_01758_),
    .Z(_01126_));
 XOR2_X1 _26895_ (.A(_01628_),
    .B(_17168_),
    .Z(_01759_));
 MUX2_X1 _26896_ (.A(_01270_),
    .B(_01759_),
    .S(_01758_),
    .Z(_01127_));
 XOR2_X1 _26897_ (.A(_01630_),
    .B(_17169_),
    .Z(_01760_));
 MUX2_X1 _26898_ (.A(_01271_),
    .B(_01760_),
    .S(_01758_),
    .Z(_01128_));
 XOR2_X2 _26899_ (.A(_17106_),
    .B(_17170_),
    .Z(_01761_));
 XOR2_X1 _26900_ (.A(_01761_),
    .B(_17138_),
    .Z(_01762_));
 XNOR2_X1 _26901_ (.A(_15642_),
    .B(_01762_),
    .ZN(_01763_));
 MUX2_X1 _26902_ (.A(_01272_),
    .B(_01763_),
    .S(_01758_),
    .Z(_01129_));
 XNOR2_X1 _26903_ (.A(_01635_),
    .B(_17171_),
    .ZN(_01764_));
 MUX2_X1 _26904_ (.A(_01273_),
    .B(_01764_),
    .S(_01758_),
    .Z(_01130_));
 XOR2_X2 _26905_ (.A(_17108_),
    .B(_17172_),
    .Z(_01765_));
 XOR2_X1 _26906_ (.A(_01765_),
    .B(_17140_),
    .Z(_01766_));
 XNOR2_X1 _26907_ (.A(_15832_),
    .B(_01766_),
    .ZN(_01767_));
 MUX2_X1 _26908_ (.A(_01275_),
    .B(_01767_),
    .S(_01758_),
    .Z(_01131_));
 XOR2_X2 _26909_ (.A(_17109_),
    .B(_17173_),
    .Z(_01768_));
 INV_X1 _26910_ (.A(_17141_),
    .ZN(_01769_));
 XNOR2_X1 _26911_ (.A(_01768_),
    .B(_01769_),
    .ZN(_01770_));
 XNOR2_X1 _26912_ (.A(_15911_),
    .B(_01770_),
    .ZN(_01771_));
 MUX2_X1 _26913_ (.A(_01276_),
    .B(_01771_),
    .S(_01758_),
    .Z(_01132_));
 MUX2_X1 _26914_ (.A(_17175_),
    .B(_01277_),
    .S(_01330_),
    .Z(_01772_));
 NAND2_X1 _26915_ (.A1(_01641_),
    .A2(_03738_),
    .ZN(_01773_));
 MUX2_X1 _26916_ (.A(_01708_),
    .B(_01772_),
    .S(_01773_),
    .Z(_01134_));
 XNOR2_X1 _26917_ (.A(_01644_),
    .B(_17176_),
    .ZN(_01774_));
 MUX2_X1 _26918_ (.A(_01278_),
    .B(_01774_),
    .S(_01758_),
    .Z(_01135_));
 XNOR2_X1 _26919_ (.A(_01647_),
    .B(_17177_),
    .ZN(_01775_));
 MUX2_X1 _26920_ (.A(_01279_),
    .B(_01775_),
    .S(_01758_),
    .Z(_01136_));
 MUX2_X1 _26921_ (.A(_17178_),
    .B(_01280_),
    .S(_01330_),
    .Z(_01776_));
 NAND2_X1 _26922_ (.A1(_01649_),
    .A2(_03738_),
    .ZN(_01777_));
 MUX2_X1 _26923_ (.A(_01727_),
    .B(_01776_),
    .S(_01777_),
    .Z(_01137_));
 XOR2_X1 _26924_ (.A(_01653_),
    .B(_17179_),
    .Z(_01778_));
 MUX2_X1 _26925_ (.A(_01281_),
    .B(_01778_),
    .S(_01758_),
    .Z(_01138_));
 XOR2_X1 _26926_ (.A(_01656_),
    .B(_17180_),
    .Z(_01779_));
 BUF_X2 _26927_ (.A(_03933_),
    .Z(_01780_));
 MUX2_X1 _26928_ (.A(_01282_),
    .B(_01779_),
    .S(_01780_),
    .Z(_01139_));
 XOR2_X1 _26929_ (.A(_01660_),
    .B(_17181_),
    .Z(_01781_));
 MUX2_X1 _26930_ (.A(_01283_),
    .B(_01781_),
    .S(_01780_),
    .Z(_01140_));
 XOR2_X1 _26931_ (.A(_01664_),
    .B(_17182_),
    .Z(_01782_));
 MUX2_X1 _26932_ (.A(_01284_),
    .B(_01782_),
    .S(_01780_),
    .Z(_01141_));
 XOR2_X1 _26933_ (.A(_01667_),
    .B(_17183_),
    .Z(_01783_));
 MUX2_X1 _26934_ (.A(_01286_),
    .B(_01783_),
    .S(_01780_),
    .Z(_01142_));
 XOR2_X1 _26935_ (.A(_01670_),
    .B(_17184_),
    .Z(_01784_));
 MUX2_X1 _26936_ (.A(_01287_),
    .B(_01784_),
    .S(_01780_),
    .Z(_01143_));
 XOR2_X1 _26937_ (.A(_01673_),
    .B(_17186_),
    .Z(_01785_));
 MUX2_X1 _26938_ (.A(_01288_),
    .B(_01785_),
    .S(_01780_),
    .Z(_01145_));
 INV_X1 _26939_ (.A(_17187_),
    .ZN(_01786_));
 XNOR2_X1 _26940_ (.A(_01676_),
    .B(_01786_),
    .ZN(_01787_));
 MUX2_X1 _26941_ (.A(_01289_),
    .B(_01787_),
    .S(_01780_),
    .Z(_01146_));
 XOR2_X1 _26942_ (.A(_17179_),
    .B(_17014_),
    .Z(_01788_));
 XNOR2_X1 _26943_ (.A(_11549_),
    .B(_13896_),
    .ZN(_01789_));
 XNOR2_X1 _26944_ (.A(_12499_),
    .B(_01033_),
    .ZN(_01790_));
 XNOR2_X1 _26945_ (.A(_01789_),
    .B(_01790_),
    .ZN(_01791_));
 MUX2_X1 _26946_ (.A(_01788_),
    .B(_01791_),
    .S(_01710_),
    .Z(_00620_));
 XOR2_X1 _26947_ (.A(_17180_),
    .B(_17015_),
    .Z(_01792_));
 INV_X1 _26948_ (.A(_01034_),
    .ZN(_01793_));
 XNOR2_X1 _26949_ (.A(_13896_),
    .B(_01793_),
    .ZN(_01794_));
 XNOR2_X1 _26950_ (.A(_01794_),
    .B(_14287_),
    .ZN(_01795_));
 XNOR2_X1 _26951_ (.A(_01690_),
    .B(_12807_),
    .ZN(_01796_));
 XNOR2_X1 _26952_ (.A(_01795_),
    .B(_01796_),
    .ZN(_01797_));
 MUX2_X1 _26953_ (.A(_01792_),
    .B(_01797_),
    .S(_01710_),
    .Z(_00621_));
 XOR2_X1 _26954_ (.A(_17181_),
    .B(_17016_),
    .Z(_01798_));
 XOR2_X1 _26955_ (.A(_12727_),
    .B(_12650_),
    .Z(_01799_));
 XNOR2_X1 _26956_ (.A(_12285_),
    .B(_01799_),
    .ZN(_01800_));
 XNOR2_X1 _26957_ (.A(_01800_),
    .B(_13017_),
    .ZN(_01801_));
 XNOR2_X1 _26958_ (.A(_01801_),
    .B(_17181_),
    .ZN(_01802_));
 MUX2_X1 _26959_ (.A(_01798_),
    .B(_01802_),
    .S(_01710_),
    .Z(_00622_));
 XOR2_X1 _26960_ (.A(_17182_),
    .B(_17017_),
    .Z(_01803_));
 XNOR2_X1 _26961_ (.A(_13287_),
    .B(_12883_),
    .ZN(_01804_));
 XNOR2_X1 _26962_ (.A(_01804_),
    .B(_13020_),
    .ZN(_01805_));
 XNOR2_X1 _26963_ (.A(_01698_),
    .B(_13094_),
    .ZN(_01806_));
 XNOR2_X1 _26964_ (.A(_01805_),
    .B(_01806_),
    .ZN(_01807_));
 XNOR2_X1 _26965_ (.A(_01807_),
    .B(_17182_),
    .ZN(_01808_));
 MUX2_X1 _26966_ (.A(_01803_),
    .B(_01808_),
    .S(_01710_),
    .Z(_00623_));
 XOR2_X1 _26967_ (.A(_17183_),
    .B(_17019_),
    .Z(_01809_));
 XNOR2_X1 _26968_ (.A(_13290_),
    .B(_01703_),
    .ZN(_01810_));
 XNOR2_X1 _26969_ (.A(_01810_),
    .B(_13216_),
    .ZN(_01811_));
 XNOR2_X1 _26970_ (.A(_01811_),
    .B(_13346_),
    .ZN(_01812_));
 XNOR2_X1 _26971_ (.A(_01812_),
    .B(_13515_),
    .ZN(_01813_));
 XNOR2_X1 _26972_ (.A(_01813_),
    .B(_17183_),
    .ZN(_01814_));
 MUX2_X1 _26973_ (.A(_01809_),
    .B(_01814_),
    .S(_01710_),
    .Z(_00624_));
 XOR2_X1 _26974_ (.A(_17184_),
    .B(_17020_),
    .Z(_01815_));
 XNOR2_X1 _26975_ (.A(_13791_),
    .B(_01035_),
    .ZN(_01816_));
 XNOR2_X1 _26976_ (.A(_13408_),
    .B(_13580_),
    .ZN(_01817_));
 XNOR2_X1 _26977_ (.A(_01816_),
    .B(_01817_),
    .ZN(_01818_));
 XOR2_X1 _26978_ (.A(_01818_),
    .B(_13217_),
    .Z(_01819_));
 MUX2_X1 _26979_ (.A(_01815_),
    .B(_01819_),
    .S(_01710_),
    .Z(_00625_));
 XOR2_X1 _26980_ (.A(_17186_),
    .B(_17021_),
    .Z(_01820_));
 XOR2_X1 _26981_ (.A(_13946_),
    .B(_01036_),
    .Z(_01821_));
 XNOR2_X1 _26982_ (.A(_01821_),
    .B(_13464_),
    .ZN(_01822_));
 XOR2_X1 _26983_ (.A(_13637_),
    .B(_13736_),
    .Z(_01823_));
 XNOR2_X1 _26984_ (.A(_01822_),
    .B(_01823_),
    .ZN(_01824_));
 BUF_X2 _26985_ (.A(_09038_),
    .Z(_01825_));
 MUX2_X1 _26986_ (.A(_01820_),
    .B(_01824_),
    .S(_01825_),
    .Z(_00626_));
 XOR2_X1 _26987_ (.A(_17187_),
    .B(_17022_),
    .Z(_01826_));
 XNOR2_X1 _26988_ (.A(_13842_),
    .B(_13895_),
    .ZN(_01827_));
 XNOR2_X1 _26989_ (.A(_13686_),
    .B(_01827_),
    .ZN(_01828_));
 XNOR2_X1 _26990_ (.A(_01828_),
    .B(_12102_),
    .ZN(_01829_));
 XNOR2_X1 _26991_ (.A(_01829_),
    .B(_01786_),
    .ZN(_01830_));
 MUX2_X1 _26992_ (.A(_01826_),
    .B(_01830_),
    .S(_01825_),
    .Z(_00627_));
 XOR2_X1 _26993_ (.A(_04132_),
    .B(_17163_),
    .Z(_01831_));
 XOR2_X1 _26994_ (.A(_01596_),
    .B(_01831_),
    .Z(_01832_));
 XNOR2_X1 _26995_ (.A(_14165_),
    .B(_01832_),
    .ZN(_01833_));
 MUX2_X1 _26996_ (.A(_01202_),
    .B(_01833_),
    .S(_01780_),
    .Z(_01154_));
 XNOR2_X1 _26997_ (.A(_09041_),
    .B(_17174_),
    .ZN(_01834_));
 XNOR2_X1 _26998_ (.A(_01599_),
    .B(_01834_),
    .ZN(_01835_));
 MUX2_X1 _26999_ (.A(_01241_),
    .B(_01835_),
    .S(_01780_),
    .Z(_01165_));
 XOR2_X1 _27000_ (.A(_17131_),
    .B(_17023_),
    .Z(_01836_));
 INV_X1 _27001_ (.A(_16694_),
    .ZN(_01837_));
 AND2_X2 _27002_ (.A1(_01837_),
    .A2(_16693_),
    .ZN(_01838_));
 INV_X1 _27003_ (.A(_16692_),
    .ZN(_01839_));
 NOR2_X1 _27004_ (.A1(_01839_),
    .A2(_16691_),
    .ZN(_01840_));
 CLKBUF_X2 _27005_ (.A(_01840_),
    .Z(_01841_));
 AND2_X1 _27006_ (.A1(_01838_),
    .A2(_01841_),
    .ZN(_01842_));
 BUF_X2 _27007_ (.A(_01842_),
    .Z(_01843_));
 NOR2_X1 _27008_ (.A1(_16689_),
    .A2(_16690_),
    .ZN(_01844_));
 CLKBUF_X2 _27009_ (.A(_01844_),
    .Z(_01845_));
 CLKBUF_X2 _27010_ (.A(_16687_),
    .Z(_01846_));
 AND2_X1 _27011_ (.A1(_01845_),
    .A2(_01846_),
    .ZN(_01847_));
 INV_X1 _27012_ (.A(_16689_),
    .ZN(_01848_));
 NOR2_X1 _27013_ (.A1(_01848_),
    .A2(_16690_),
    .ZN(_01849_));
 BUF_X1 _27014_ (.A(_01849_),
    .Z(_01850_));
 CLKBUF_X2 _27015_ (.A(_01850_),
    .Z(_01851_));
 BUF_X2 _27016_ (.A(_01851_),
    .Z(_01852_));
 OAI21_X1 _27017_ (.A(_01843_),
    .B1(_01847_),
    .B2(_01852_),
    .ZN(_01853_));
 AND2_X1 _27018_ (.A1(_01839_),
    .A2(_16691_),
    .ZN(_01854_));
 AND2_X1 _27019_ (.A1(_01838_),
    .A2(_01854_),
    .ZN(_01855_));
 AND2_X2 _27020_ (.A1(_16688_),
    .A2(_16687_),
    .ZN(_01856_));
 AND2_X1 _27021_ (.A1(_01856_),
    .A2(_01844_),
    .ZN(_01857_));
 BUF_X2 _27022_ (.A(_01857_),
    .Z(_01858_));
 NAND2_X1 _27023_ (.A1(_01855_),
    .A2(_01858_),
    .ZN(_01859_));
 INV_X1 _27024_ (.A(_16688_),
    .ZN(_01860_));
 CLKBUF_X2 _27025_ (.A(_01860_),
    .Z(_01861_));
 AND2_X1 _27026_ (.A1(_01844_),
    .A2(_01861_),
    .ZN(_01862_));
 NAND3_X1 _27027_ (.A1(_01862_),
    .A2(_01838_),
    .A3(_01854_),
    .ZN(_01863_));
 NAND2_X1 _27028_ (.A1(_01859_),
    .A2(_01863_),
    .ZN(_01864_));
 INV_X1 _27029_ (.A(_16690_),
    .ZN(_01865_));
 NOR2_X1 _27030_ (.A1(_01865_),
    .A2(_16689_),
    .ZN(_01866_));
 CLKBUF_X2 _27031_ (.A(_01866_),
    .Z(_01867_));
 AND2_X1 _27032_ (.A1(_01867_),
    .A2(_16687_),
    .ZN(_01868_));
 AND2_X1 _27033_ (.A1(_16689_),
    .A2(_16690_),
    .ZN(_01869_));
 AND2_X2 _27034_ (.A1(_01869_),
    .A2(_01856_),
    .ZN(_01870_));
 OAI21_X1 _27035_ (.A(_01855_),
    .B1(_01868_),
    .B2(_01870_),
    .ZN(_01871_));
 NOR2_X2 _27036_ (.A1(_16688_),
    .A2(_16687_),
    .ZN(_01872_));
 AND2_X1 _27037_ (.A1(_01850_),
    .A2(_01872_),
    .ZN(_01873_));
 NOR2_X1 _27038_ (.A1(_16692_),
    .A2(_16691_),
    .ZN(_01874_));
 CLKBUF_X2 _27039_ (.A(_01874_),
    .Z(_01875_));
 NAND3_X1 _27040_ (.A1(_01873_),
    .A2(_01838_),
    .A3(_01875_),
    .ZN(_01876_));
 INV_X1 _27041_ (.A(_01862_),
    .ZN(_01877_));
 AND2_X1 _27042_ (.A1(_01838_),
    .A2(_01874_),
    .ZN(_01878_));
 INV_X1 _27043_ (.A(_01878_),
    .ZN(_01879_));
 OAI211_X1 _27044_ (.A(_01871_),
    .B(_01876_),
    .C1(_01877_),
    .C2(_01879_),
    .ZN(_01880_));
 NOR2_X2 _27045_ (.A1(_01860_),
    .A2(_16687_),
    .ZN(_01881_));
 NOR3_X1 _27046_ (.A1(_01881_),
    .A2(_16689_),
    .A3(_01865_),
    .ZN(_01882_));
 AOI211_X1 _27047_ (.A(_01864_),
    .B(_01880_),
    .C1(_01843_),
    .C2(_01882_),
    .ZN(_01883_));
 AND2_X1 _27048_ (.A1(_01850_),
    .A2(_16687_),
    .ZN(_01884_));
 BUF_X2 _27049_ (.A(_01838_),
    .Z(_01885_));
 AND2_X2 _27050_ (.A1(_16692_),
    .A2(_16691_),
    .ZN(_01886_));
 BUF_X2 _27051_ (.A(_01886_),
    .Z(_01887_));
 NAND3_X1 _27052_ (.A1(_01884_),
    .A2(_01885_),
    .A3(_01887_),
    .ZN(_01888_));
 AND2_X1 _27053_ (.A1(_01838_),
    .A2(_01886_),
    .ZN(_01889_));
 BUF_X2 _27054_ (.A(_01889_),
    .Z(_01890_));
 NAND2_X1 _27055_ (.A1(_01890_),
    .A2(_01858_),
    .ZN(_01891_));
 AND2_X1 _27056_ (.A1(_01888_),
    .A2(_01891_),
    .ZN(_01892_));
 INV_X1 _27057_ (.A(_01851_),
    .ZN(_01893_));
 CLKBUF_X2 _27058_ (.A(_01881_),
    .Z(_01894_));
 NOR2_X1 _27059_ (.A1(_01893_),
    .A2(_01894_),
    .ZN(_01895_));
 NOR2_X2 _27060_ (.A1(_01837_),
    .A2(_16693_),
    .ZN(_01896_));
 AND2_X1 _27061_ (.A1(_01896_),
    .A2(_01874_),
    .ZN(_01897_));
 BUF_X2 _27062_ (.A(_01897_),
    .Z(_01898_));
 NAND2_X1 _27063_ (.A1(_01895_),
    .A2(_01898_),
    .ZN(_01899_));
 AND4_X1 _27064_ (.A1(_01853_),
    .A2(_01883_),
    .A3(_01892_),
    .A4(_01899_),
    .ZN(_01900_));
 AND2_X2 _27065_ (.A1(_01896_),
    .A2(_01840_),
    .ZN(_01901_));
 AND2_X1 _27066_ (.A1(_01869_),
    .A2(_01861_),
    .ZN(_01902_));
 CLKBUF_X2 _27067_ (.A(_01902_),
    .Z(_01903_));
 OAI21_X1 _27068_ (.A(_01901_),
    .B1(_01870_),
    .B2(_01903_),
    .ZN(_01904_));
 BUF_X2 _27069_ (.A(_01867_),
    .Z(_01905_));
 INV_X1 _27070_ (.A(_16687_),
    .ZN(_01906_));
 NOR2_X2 _27071_ (.A1(_01906_),
    .A2(_16688_),
    .ZN(_01907_));
 NAND4_X1 _27072_ (.A1(_01905_),
    .A2(_01907_),
    .A3(_01896_),
    .A4(_01841_),
    .ZN(_01908_));
 AND2_X1 _27073_ (.A1(_01904_),
    .A2(_01908_),
    .ZN(_01909_));
 AND2_X1 _27074_ (.A1(_01881_),
    .A2(_01869_),
    .ZN(_01910_));
 BUF_X2 _27075_ (.A(_01910_),
    .Z(_01911_));
 AND2_X1 _27076_ (.A1(_01907_),
    .A2(_01869_),
    .ZN(_01912_));
 OAI21_X1 _27077_ (.A(_01890_),
    .B1(_01911_),
    .B2(_01912_),
    .ZN(_01913_));
 AND2_X1 _27078_ (.A1(_01866_),
    .A2(_01856_),
    .ZN(_01914_));
 BUF_X2 _27079_ (.A(_01914_),
    .Z(_01915_));
 NAND3_X1 _27080_ (.A1(_01915_),
    .A2(_01885_),
    .A3(_01886_),
    .ZN(_01916_));
 NAND2_X1 _27081_ (.A1(_01913_),
    .A2(_01916_),
    .ZN(_01917_));
 INV_X1 _27082_ (.A(_01917_),
    .ZN(_01918_));
 INV_X1 _27083_ (.A(_01867_),
    .ZN(_01919_));
 CLKBUF_X2 _27084_ (.A(_01906_),
    .Z(_01920_));
 INV_X1 _27085_ (.A(_01869_),
    .ZN(_01921_));
 CLKBUF_X2 _27086_ (.A(_01872_),
    .Z(_01922_));
 OAI22_X1 _27087_ (.A1(_01919_),
    .A2(_01920_),
    .B1(_01921_),
    .B2(_01922_),
    .ZN(_01923_));
 AND2_X1 _27088_ (.A1(_01845_),
    .A2(_01906_),
    .ZN(_01924_));
 OAI21_X1 _27089_ (.A(_01898_),
    .B1(_01923_),
    .B2(_01924_),
    .ZN(_01925_));
 AND2_X1 _27090_ (.A1(_01896_),
    .A2(_01886_),
    .ZN(_01926_));
 INV_X2 _27091_ (.A(_01845_),
    .ZN(_01927_));
 NOR2_X1 _27092_ (.A1(_01927_),
    .A2(_01907_),
    .ZN(_01928_));
 AND2_X1 _27093_ (.A1(_01926_),
    .A2(_01928_),
    .ZN(_01929_));
 INV_X1 _27094_ (.A(_01929_),
    .ZN(_01930_));
 AND4_X1 _27095_ (.A1(_01909_),
    .A2(_01918_),
    .A3(_01925_),
    .A4(_01930_),
    .ZN(_01931_));
 NOR2_X2 _27096_ (.A1(_16694_),
    .A2(_16693_),
    .ZN(_01932_));
 AND2_X1 _27097_ (.A1(_01841_),
    .A2(_01932_),
    .ZN(_01933_));
 BUF_X2 _27098_ (.A(_01933_),
    .Z(_01934_));
 NOR3_X2 _27099_ (.A1(_01872_),
    .A2(_01848_),
    .A3(_16690_),
    .ZN(_01935_));
 INV_X1 _27100_ (.A(_01856_),
    .ZN(_01936_));
 AND2_X1 _27101_ (.A1(_01935_),
    .A2(_01936_),
    .ZN(_01937_));
 CLKBUF_X2 _27102_ (.A(_01869_),
    .Z(_01938_));
 AND2_X1 _27103_ (.A1(_01938_),
    .A2(_01920_),
    .ZN(_01939_));
 OAI21_X1 _27104_ (.A(_01934_),
    .B1(_01937_),
    .B2(_01939_),
    .ZN(_01940_));
 AND2_X1 _27105_ (.A1(_16694_),
    .A2(_16693_),
    .ZN(_01941_));
 AND2_X1 _27106_ (.A1(_01840_),
    .A2(_01941_),
    .ZN(_01942_));
 BUF_X2 _27107_ (.A(_01942_),
    .Z(_01943_));
 INV_X1 _27108_ (.A(_01858_),
    .ZN(_01944_));
 AND2_X2 _27109_ (.A1(_01872_),
    .A2(_01845_),
    .ZN(_01945_));
 INV_X1 _27110_ (.A(_01945_),
    .ZN(_01946_));
 NAND2_X1 _27111_ (.A1(_01944_),
    .A2(_01946_),
    .ZN(_01947_));
 AND2_X1 _27112_ (.A1(_01850_),
    .A2(_01861_),
    .ZN(_01948_));
 BUF_X2 _27113_ (.A(_01948_),
    .Z(_01949_));
 OAI21_X1 _27114_ (.A(_01943_),
    .B1(_01947_),
    .B2(_01949_),
    .ZN(_01950_));
 AND2_X1 _27115_ (.A1(_01854_),
    .A2(_01932_),
    .ZN(_01951_));
 BUF_X2 _27116_ (.A(_01951_),
    .Z(_01952_));
 AND2_X2 _27117_ (.A1(_01845_),
    .A2(_16688_),
    .ZN(_01953_));
 CLKBUF_X2 _27118_ (.A(_16688_),
    .Z(_01954_));
 AND2_X1 _27119_ (.A1(_01850_),
    .A2(_01954_),
    .ZN(_01955_));
 BUF_X2 _27120_ (.A(_01955_),
    .Z(_01956_));
 AND2_X1 _27121_ (.A1(_01932_),
    .A2(_01874_),
    .ZN(_01957_));
 CLKBUF_X2 _27122_ (.A(_01957_),
    .Z(_01958_));
 AOI22_X1 _27123_ (.A1(_01952_),
    .A2(_01953_),
    .B1(_01956_),
    .B2(_01958_),
    .ZN(_01959_));
 AND2_X1 _27124_ (.A1(_01854_),
    .A2(_01896_),
    .ZN(_01960_));
 BUF_X2 _27125_ (.A(_01960_),
    .Z(_01961_));
 NOR3_X1 _27126_ (.A1(_01927_),
    .A2(_01856_),
    .A3(_01922_),
    .ZN(_01962_));
 AND2_X2 _27127_ (.A1(_01869_),
    .A2(_01954_),
    .ZN(_01963_));
 OAI21_X1 _27128_ (.A(_01961_),
    .B1(_01962_),
    .B2(_01963_),
    .ZN(_01964_));
 AND4_X1 _27129_ (.A1(_01940_),
    .A2(_01950_),
    .A3(_01959_),
    .A4(_01964_),
    .ZN(_01965_));
 NAND2_X1 _27130_ (.A1(_01842_),
    .A2(_01911_),
    .ZN(_01966_));
 NAND2_X1 _27131_ (.A1(_01933_),
    .A2(_01870_),
    .ZN(_01967_));
 AND2_X2 _27132_ (.A1(_01867_),
    .A2(_01907_),
    .ZN(_01968_));
 INV_X1 _27133_ (.A(_01968_),
    .ZN(_01969_));
 AND2_X1 _27134_ (.A1(_01941_),
    .A2(_01874_),
    .ZN(_01970_));
 INV_X1 _27135_ (.A(_01970_),
    .ZN(_01971_));
 OAI211_X1 _27136_ (.A(_01966_),
    .B(_01967_),
    .C1(_01969_),
    .C2(_01971_),
    .ZN(_01972_));
 CLKBUF_X2 _27137_ (.A(_01901_),
    .Z(_01973_));
 AND2_X1 _27138_ (.A1(_01886_),
    .A2(_01932_),
    .ZN(_01974_));
 BUF_X2 _27139_ (.A(_01974_),
    .Z(_01975_));
 AOI22_X1 _27140_ (.A1(_01973_),
    .A2(_01873_),
    .B1(_01870_),
    .B2(_01975_),
    .ZN(_01976_));
 NAND2_X1 _27141_ (.A1(_01958_),
    .A2(_01953_),
    .ZN(_01977_));
 AND2_X1 _27142_ (.A1(_01869_),
    .A2(_01872_),
    .ZN(_01978_));
 BUF_X2 _27143_ (.A(_01978_),
    .Z(_01979_));
 CLKBUF_X2 _27144_ (.A(_01896_),
    .Z(_01980_));
 NAND3_X1 _27145_ (.A1(_01979_),
    .A2(_01980_),
    .A3(_01887_),
    .ZN(_01981_));
 NAND3_X1 _27146_ (.A1(_01976_),
    .A2(_01977_),
    .A3(_01981_),
    .ZN(_01982_));
 BUF_X2 _27147_ (.A(_01926_),
    .Z(_01983_));
 AOI211_X1 _27148_ (.A(_01972_),
    .B(_01982_),
    .C1(_01983_),
    .C2(_01895_),
    .ZN(_01984_));
 AND4_X1 _27149_ (.A1(_01900_),
    .A2(_01931_),
    .A3(_01965_),
    .A4(_01984_),
    .ZN(_01985_));
 NOR2_X1 _27150_ (.A1(_01910_),
    .A2(_01912_),
    .ZN(_01986_));
 AND2_X1 _27151_ (.A1(_01907_),
    .A2(_01850_),
    .ZN(_01987_));
 INV_X1 _27152_ (.A(_01987_),
    .ZN(_01988_));
 AND2_X1 _27153_ (.A1(_01866_),
    .A2(_16688_),
    .ZN(_01989_));
 INV_X1 _27154_ (.A(_01989_),
    .ZN(_01990_));
 NAND4_X1 _27155_ (.A1(_01986_),
    .A2(_01969_),
    .A3(_01988_),
    .A4(_01990_),
    .ZN(_01991_));
 BUF_X2 _27156_ (.A(_01957_),
    .Z(_01992_));
 NAND2_X1 _27157_ (.A1(_01991_),
    .A2(_01992_),
    .ZN(_01993_));
 NOR3_X1 _27158_ (.A1(_01907_),
    .A2(_16689_),
    .A3(_01865_),
    .ZN(_01994_));
 INV_X1 _27159_ (.A(_01881_),
    .ZN(_01995_));
 AND2_X1 _27160_ (.A1(_01994_),
    .A2(_01995_),
    .ZN(_01996_));
 OAI21_X1 _27161_ (.A(_01951_),
    .B1(_01996_),
    .B2(_01937_),
    .ZN(_01997_));
 NAND2_X1 _27162_ (.A1(_01975_),
    .A2(_01903_),
    .ZN(_01998_));
 AND2_X1 _27163_ (.A1(_01881_),
    .A2(_01850_),
    .ZN(_01999_));
 BUF_X2 _27164_ (.A(_01999_),
    .Z(_02000_));
 AND2_X1 _27165_ (.A1(_01867_),
    .A2(_01922_),
    .ZN(_02001_));
 OAI21_X1 _27166_ (.A(_01975_),
    .B1(_02000_),
    .B2(_02001_),
    .ZN(_02002_));
 AND3_X1 _27167_ (.A1(_01997_),
    .A2(_01998_),
    .A3(_02002_),
    .ZN(_02003_));
 AND2_X1 _27168_ (.A1(_01994_),
    .A2(_01942_),
    .ZN(_02004_));
 INV_X1 _27169_ (.A(_01872_),
    .ZN(_02005_));
 AND2_X1 _27170_ (.A1(_02005_),
    .A2(_01866_),
    .ZN(_02006_));
 NOR2_X1 _27171_ (.A1(_01927_),
    .A2(_01872_),
    .ZN(_02007_));
 AOI221_X1 _27172_ (.A(_02004_),
    .B1(_02006_),
    .B2(_01933_),
    .C1(_01975_),
    .C2(_02007_),
    .ZN(_02008_));
 CLKBUF_X2 _27173_ (.A(_01936_),
    .Z(_02009_));
 AND3_X1 _27174_ (.A1(_02009_),
    .A2(_01941_),
    .A3(_01874_),
    .ZN(_02010_));
 OAI21_X1 _27175_ (.A(_02010_),
    .B1(_01938_),
    .B2(_01953_),
    .ZN(_02011_));
 BUF_X2 _27176_ (.A(_01862_),
    .Z(_02012_));
 NAND3_X1 _27177_ (.A1(_02012_),
    .A2(_01885_),
    .A3(_01886_),
    .ZN(_02013_));
 BUF_X2 _27178_ (.A(_01855_),
    .Z(_02014_));
 NAND2_X1 _27179_ (.A1(_02014_),
    .A2(_01956_),
    .ZN(_02015_));
 AND3_X1 _27180_ (.A1(_02011_),
    .A2(_02013_),
    .A3(_02015_),
    .ZN(_02016_));
 AND2_X1 _27181_ (.A1(_01886_),
    .A2(_01941_),
    .ZN(_02017_));
 BUF_X2 _27182_ (.A(_02017_),
    .Z(_02018_));
 INV_X1 _27183_ (.A(_02018_),
    .ZN(_02019_));
 INV_X1 _27184_ (.A(_01910_),
    .ZN(_02020_));
 INV_X1 _27185_ (.A(_01873_),
    .ZN(_02021_));
 AOI21_X1 _27186_ (.A(_02019_),
    .B1(_02020_),
    .B2(_02021_),
    .ZN(_02022_));
 AND2_X1 _27187_ (.A1(_01914_),
    .A2(_01970_),
    .ZN(_02023_));
 AND2_X1 _27188_ (.A1(_01907_),
    .A2(_01845_),
    .ZN(_02024_));
 AND2_X1 _27189_ (.A1(_02024_),
    .A2(_02017_),
    .ZN(_02025_));
 NOR2_X1 _27190_ (.A1(_01927_),
    .A2(_01856_),
    .ZN(_02026_));
 AND2_X1 _27191_ (.A1(_01933_),
    .A2(_02026_),
    .ZN(_02027_));
 NOR4_X1 _27192_ (.A1(_02022_),
    .A2(_02023_),
    .A3(_02025_),
    .A4(_02027_),
    .ZN(_02028_));
 AND4_X1 _27193_ (.A1(_02003_),
    .A2(_02008_),
    .A3(_02016_),
    .A4(_02028_),
    .ZN(_02029_));
 AND2_X1 _27194_ (.A1(_01854_),
    .A2(_01941_),
    .ZN(_02030_));
 BUF_X2 _27195_ (.A(_02030_),
    .Z(_02031_));
 BUF_X2 _27196_ (.A(_01987_),
    .Z(_02032_));
 AND2_X1 _27197_ (.A1(_01881_),
    .A2(_01844_),
    .ZN(_02033_));
 OAI21_X1 _27198_ (.A(_02031_),
    .B1(_02032_),
    .B2(_02033_),
    .ZN(_02034_));
 BUF_X2 _27199_ (.A(_01989_),
    .Z(_02035_));
 AND2_X1 _27200_ (.A1(_01866_),
    .A2(_01861_),
    .ZN(_02036_));
 BUF_X2 _27201_ (.A(_02036_),
    .Z(_02037_));
 OAI21_X1 _27202_ (.A(_02031_),
    .B1(_02035_),
    .B2(_02037_),
    .ZN(_02038_));
 AND2_X1 _27203_ (.A1(_01938_),
    .A2(_01846_),
    .ZN(_02039_));
 AOI21_X1 _27204_ (.A(_16689_),
    .B1(_01861_),
    .B2(_01865_),
    .ZN(_02040_));
 AOI22_X1 _27205_ (.A1(_01943_),
    .A2(_02039_),
    .B1(_02018_),
    .B2(_02040_),
    .ZN(_02041_));
 BUF_X2 _27206_ (.A(_01912_),
    .Z(_02042_));
 OAI21_X1 _27207_ (.A(_02031_),
    .B1(_01911_),
    .B2(_02042_),
    .ZN(_02043_));
 AND4_X1 _27208_ (.A1(_02034_),
    .A2(_02038_),
    .A3(_02041_),
    .A4(_02043_),
    .ZN(_02044_));
 AND2_X1 _27209_ (.A1(_01945_),
    .A2(_01992_),
    .ZN(_02045_));
 OR3_X1 _27210_ (.A1(_01868_),
    .A2(_01939_),
    .A3(_01903_),
    .ZN(_02046_));
 BUF_X2 _27211_ (.A(_01878_),
    .Z(_02047_));
 AOI21_X1 _27212_ (.A(_02045_),
    .B1(_02046_),
    .B2(_02047_),
    .ZN(_02048_));
 AND4_X1 _27213_ (.A1(_01993_),
    .A2(_02029_),
    .A3(_02044_),
    .A4(_02048_),
    .ZN(_02049_));
 AND2_X1 _27214_ (.A1(_01985_),
    .A2(_02049_),
    .ZN(_02050_));
 AND2_X1 _27215_ (.A1(_02036_),
    .A2(_01970_),
    .ZN(_02051_));
 INV_X1 _27216_ (.A(_02051_),
    .ZN(_02052_));
 AND2_X1 _27217_ (.A1(_02030_),
    .A2(_01914_),
    .ZN(_02053_));
 AND2_X1 _27218_ (.A1(_02030_),
    .A2(_02000_),
    .ZN(_02054_));
 AND3_X1 _27219_ (.A1(_02033_),
    .A2(_01854_),
    .A3(_01941_),
    .ZN(_02055_));
 OR2_X1 _27220_ (.A1(_02054_),
    .A2(_02055_),
    .ZN(_02056_));
 NOR2_X2 _27221_ (.A1(_01921_),
    .A2(_01881_),
    .ZN(_02057_));
 AOI211_X1 _27222_ (.A(_02053_),
    .B(_02056_),
    .C1(_02057_),
    .C2(_02031_),
    .ZN(_02058_));
 BUF_X2 _27223_ (.A(_01970_),
    .Z(_02059_));
 OAI21_X1 _27224_ (.A(_02059_),
    .B1(_01935_),
    .B2(_01945_),
    .ZN(_02060_));
 CLKBUF_X2 _27225_ (.A(_01938_),
    .Z(_02061_));
 OAI211_X1 _27226_ (.A(_02059_),
    .B(_02061_),
    .C1(_01954_),
    .C2(_01846_),
    .ZN(_02062_));
 AND4_X1 _27227_ (.A1(_02052_),
    .A2(_02058_),
    .A3(_02060_),
    .A4(_02062_),
    .ZN(_02063_));
 OAI21_X1 _27228_ (.A(_02018_),
    .B1(_01968_),
    .B2(_01939_),
    .ZN(_02064_));
 INV_X1 _27229_ (.A(_01943_),
    .ZN(_02065_));
 INV_X1 _27230_ (.A(_02033_),
    .ZN(_02066_));
 AOI21_X1 _27231_ (.A(_02065_),
    .B1(_02066_),
    .B2(_01877_),
    .ZN(_02067_));
 INV_X1 _27232_ (.A(_01955_),
    .ZN(_02068_));
 AOI21_X1 _27233_ (.A(_02065_),
    .B1(_01988_),
    .B2(_02068_),
    .ZN(_02069_));
 NOR2_X1 _27234_ (.A1(_02067_),
    .A2(_02069_),
    .ZN(_02070_));
 OAI21_X1 _27235_ (.A(_02018_),
    .B1(_01949_),
    .B2(_02026_),
    .ZN(_02071_));
 INV_X1 _27236_ (.A(_01907_),
    .ZN(_02072_));
 OAI211_X1 _27237_ (.A(_02072_),
    .B(_01943_),
    .C1(_02057_),
    .C2(_01905_),
    .ZN(_02073_));
 AND4_X1 _27238_ (.A1(_02064_),
    .A2(_02070_),
    .A3(_02071_),
    .A4(_02073_),
    .ZN(_02074_));
 OAI21_X1 _27239_ (.A(_01961_),
    .B1(_01956_),
    .B2(_01847_),
    .ZN(_02075_));
 AND2_X1 _27240_ (.A1(_02006_),
    .A2(_02009_),
    .ZN(_02076_));
 INV_X1 _27241_ (.A(_01870_),
    .ZN(_02077_));
 INV_X1 _27242_ (.A(_01979_),
    .ZN(_02078_));
 NAND2_X1 _27243_ (.A1(_02077_),
    .A2(_02078_),
    .ZN(_02079_));
 OAI21_X1 _27244_ (.A(_01960_),
    .B1(_02076_),
    .B2(_02079_),
    .ZN(_02080_));
 NAND2_X1 _27245_ (.A1(_01898_),
    .A2(_02037_),
    .ZN(_02081_));
 OAI21_X1 _27246_ (.A(_01897_),
    .B1(_01947_),
    .B2(_02032_),
    .ZN(_02082_));
 AND4_X1 _27247_ (.A1(_02075_),
    .A2(_02080_),
    .A3(_02081_),
    .A4(_02082_),
    .ZN(_02083_));
 NAND2_X1 _27248_ (.A1(_01989_),
    .A2(_01926_),
    .ZN(_02084_));
 NAND2_X1 _27249_ (.A1(_01911_),
    .A2(_01926_),
    .ZN(_02085_));
 AND2_X1 _27250_ (.A1(_02084_),
    .A2(_02085_),
    .ZN(_02086_));
 NAND2_X1 _27251_ (.A1(_01901_),
    .A2(_01945_),
    .ZN(_02087_));
 BUF_X2 _27252_ (.A(_01861_),
    .Z(_02088_));
 OAI221_X1 _27253_ (.A(_01973_),
    .B1(_02088_),
    .B2(_01920_),
    .C1(_02061_),
    .C2(_01905_),
    .ZN(_02089_));
 OAI21_X1 _27254_ (.A(_01983_),
    .B1(_01895_),
    .B2(_02012_),
    .ZN(_02090_));
 AND4_X1 _27255_ (.A1(_02086_),
    .A2(_02087_),
    .A3(_02089_),
    .A4(_02090_),
    .ZN(_02091_));
 NAND4_X2 _27256_ (.A1(_02063_),
    .A2(_02074_),
    .A3(_02083_),
    .A4(_02091_),
    .ZN(_02092_));
 OAI21_X1 _27257_ (.A(_02014_),
    .B1(_02076_),
    .B2(_01870_),
    .ZN(_02093_));
 CLKBUF_X2 _27258_ (.A(_01854_),
    .Z(_02094_));
 NAND4_X1 _27259_ (.A1(_01885_),
    .A2(_02094_),
    .A3(_01846_),
    .A4(_01845_),
    .ZN(_02095_));
 OAI21_X1 _27260_ (.A(_02014_),
    .B1(_02032_),
    .B2(_02000_),
    .ZN(_02096_));
 AND3_X1 _27261_ (.A1(_02093_),
    .A2(_02095_),
    .A3(_02096_),
    .ZN(_02097_));
 AND2_X1 _27262_ (.A1(_01849_),
    .A2(_01856_),
    .ZN(_02098_));
 AND2_X1 _27263_ (.A1(_01842_),
    .A2(_02098_),
    .ZN(_02099_));
 INV_X1 _27264_ (.A(_01842_),
    .ZN(_02100_));
 INV_X1 _27265_ (.A(_01963_),
    .ZN(_02101_));
 AOI21_X1 _27266_ (.A(_02100_),
    .B1(_01969_),
    .B2(_02101_),
    .ZN(_02102_));
 CLKBUF_X2 _27267_ (.A(_01845_),
    .Z(_02103_));
 AOI211_X1 _27268_ (.A(_02099_),
    .B(_02102_),
    .C1(_02103_),
    .C2(_01842_),
    .ZN(_02104_));
 INV_X1 _27269_ (.A(_02039_),
    .ZN(_02105_));
 AOI21_X1 _27270_ (.A(_01879_),
    .B1(_01990_),
    .B2(_02105_),
    .ZN(_02106_));
 INV_X1 _27271_ (.A(_02098_),
    .ZN(_02107_));
 BUF_X2 _27272_ (.A(_02024_),
    .Z(_02108_));
 INV_X1 _27273_ (.A(_02108_),
    .ZN(_02109_));
 NAND2_X1 _27274_ (.A1(_02107_),
    .A2(_02109_),
    .ZN(_02110_));
 AOI21_X1 _27275_ (.A(_02106_),
    .B1(_02047_),
    .B2(_02110_),
    .ZN(_02111_));
 NAND2_X1 _27276_ (.A1(_01889_),
    .A2(_01847_),
    .ZN(_02112_));
 AND2_X2 _27277_ (.A1(_01867_),
    .A2(_01881_),
    .ZN(_02113_));
 OAI21_X1 _27278_ (.A(_01889_),
    .B1(_02113_),
    .B2(_02036_),
    .ZN(_02114_));
 OAI21_X1 _27279_ (.A(_01889_),
    .B1(_02098_),
    .B2(_01948_),
    .ZN(_02115_));
 OAI21_X1 _27280_ (.A(_01889_),
    .B1(_01912_),
    .B2(_01963_),
    .ZN(_02116_));
 AND4_X1 _27281_ (.A1(_02112_),
    .A2(_02114_),
    .A3(_02115_),
    .A4(_02116_),
    .ZN(_02117_));
 AND4_X1 _27282_ (.A1(_02097_),
    .A2(_02104_),
    .A3(_02111_),
    .A4(_02117_),
    .ZN(_02118_));
 AND3_X1 _27283_ (.A1(_01958_),
    .A2(_01938_),
    .A3(_01894_),
    .ZN(_02119_));
 AND4_X1 _27284_ (.A1(_01995_),
    .A2(_01958_),
    .A3(_02072_),
    .A4(_01851_),
    .ZN(_02120_));
 AOI211_X1 _27285_ (.A(_02119_),
    .B(_02120_),
    .C1(_01903_),
    .C2(_01992_),
    .ZN(_02121_));
 NAND2_X1 _27286_ (.A1(_02107_),
    .A2(_02021_),
    .ZN(_02122_));
 AND2_X1 _27287_ (.A1(_02122_),
    .A2(_01952_),
    .ZN(_02123_));
 NAND2_X1 _27288_ (.A1(_01951_),
    .A2(_02012_),
    .ZN(_02124_));
 INV_X2 _27289_ (.A(_01951_),
    .ZN(_02125_));
 OAI21_X1 _27290_ (.A(_02124_),
    .B1(_02125_),
    .B2(_02066_),
    .ZN(_02126_));
 NAND2_X1 _27291_ (.A1(_01951_),
    .A2(_02037_),
    .ZN(_02127_));
 OAI21_X1 _27292_ (.A(_02127_),
    .B1(_02125_),
    .B2(_01990_),
    .ZN(_02128_));
 NAND2_X1 _27293_ (.A1(_01952_),
    .A2(_01903_),
    .ZN(_02129_));
 OAI21_X1 _27294_ (.A(_02129_),
    .B1(_02125_),
    .B2(_02077_),
    .ZN(_02130_));
 NOR4_X1 _27295_ (.A1(_02123_),
    .A2(_02126_),
    .A3(_02128_),
    .A4(_02130_),
    .ZN(_02131_));
 BUF_X2 _27296_ (.A(_01975_),
    .Z(_02132_));
 OAI21_X1 _27297_ (.A(_02132_),
    .B1(_01989_),
    .B2(_01939_),
    .ZN(_02133_));
 OAI21_X1 _27298_ (.A(_01934_),
    .B1(_02006_),
    .B2(_02042_),
    .ZN(_02134_));
 OAI21_X1 _27299_ (.A(_01933_),
    .B1(_01956_),
    .B2(_02026_),
    .ZN(_02135_));
 OAI211_X1 _27300_ (.A(_01975_),
    .B(_01846_),
    .C1(_02103_),
    .C2(_01851_),
    .ZN(_02136_));
 AND4_X1 _27301_ (.A1(_02133_),
    .A2(_02134_),
    .A3(_02135_),
    .A4(_02136_),
    .ZN(_02137_));
 NAND4_X2 _27302_ (.A1(_02118_),
    .A2(_02121_),
    .A3(_02131_),
    .A4(_02137_),
    .ZN(_02138_));
 NOR2_X4 _27303_ (.A1(_02092_),
    .A2(_02138_),
    .ZN(_02139_));
 XNOR2_X2 _27304_ (.A(_02050_),
    .B(_02139_),
    .ZN(_02140_));
 INV_X1 _27305_ (.A(_02140_),
    .ZN(_02141_));
 AND2_X1 _27306_ (.A1(_16769_),
    .A2(_16770_),
    .ZN(_02142_));
 INV_X1 _27307_ (.A(_02142_),
    .ZN(_02143_));
 NOR2_X1 _27308_ (.A1(_16768_),
    .A2(_16767_),
    .ZN(_02144_));
 BUF_X2 _27309_ (.A(_02144_),
    .Z(_02145_));
 NOR2_X1 _27310_ (.A1(_02143_),
    .A2(_02145_),
    .ZN(_02146_));
 INV_X1 _27311_ (.A(_16774_),
    .ZN(_02147_));
 NOR2_X1 _27312_ (.A1(_02147_),
    .A2(_16773_),
    .ZN(_02148_));
 NOR2_X1 _27313_ (.A1(_16772_),
    .A2(_16771_),
    .ZN(_02149_));
 CLKBUF_X2 _27314_ (.A(_02149_),
    .Z(_02150_));
 AND2_X1 _27315_ (.A1(_02148_),
    .A2(_02150_),
    .ZN(_02151_));
 BUF_X2 _27316_ (.A(_02151_),
    .Z(_02152_));
 AND2_X1 _27317_ (.A1(_02146_),
    .A2(_02152_),
    .ZN(_02153_));
 INV_X1 _27318_ (.A(_02153_),
    .ZN(_02154_));
 INV_X1 _27319_ (.A(_16770_),
    .ZN(_02155_));
 NOR2_X1 _27320_ (.A1(_02155_),
    .A2(_16769_),
    .ZN(_02156_));
 CLKBUF_X2 _27321_ (.A(_02156_),
    .Z(_02157_));
 BUF_X2 _27322_ (.A(_16767_),
    .Z(_02158_));
 AND2_X1 _27323_ (.A1(_02157_),
    .A2(_02158_),
    .ZN(_02159_));
 NOR2_X1 _27324_ (.A1(_16769_),
    .A2(_16770_),
    .ZN(_02160_));
 CLKBUF_X2 _27325_ (.A(_02160_),
    .Z(_02161_));
 CLKBUF_X2 _27326_ (.A(_02161_),
    .Z(_02162_));
 INV_X1 _27327_ (.A(_02158_),
    .ZN(_02163_));
 AND2_X1 _27328_ (.A1(_02162_),
    .A2(_02163_),
    .ZN(_02164_));
 OAI21_X1 _27329_ (.A(_02151_),
    .B1(_02159_),
    .B2(_02164_),
    .ZN(_02165_));
 AND2_X2 _27330_ (.A1(_16768_),
    .A2(_02158_),
    .ZN(_02166_));
 AND2_X1 _27331_ (.A1(_02142_),
    .A2(_02166_),
    .ZN(_02167_));
 AND2_X1 _27332_ (.A1(_02147_),
    .A2(_16773_),
    .ZN(_02168_));
 INV_X1 _27333_ (.A(_16772_),
    .ZN(_02169_));
 AND2_X1 _27334_ (.A1(_02169_),
    .A2(_16771_),
    .ZN(_02170_));
 CLKBUF_X2 _27335_ (.A(_02170_),
    .Z(_02171_));
 AND3_X1 _27336_ (.A1(_02167_),
    .A2(_02168_),
    .A3(_02171_),
    .ZN(_02172_));
 AND2_X1 _27337_ (.A1(_02170_),
    .A2(_02168_),
    .ZN(_02173_));
 INV_X1 _27338_ (.A(_02145_),
    .ZN(_02174_));
 NAND2_X1 _27339_ (.A1(_02174_),
    .A2(_02161_),
    .ZN(_02175_));
 INV_X1 _27340_ (.A(_02175_),
    .ZN(_02176_));
 AND2_X1 _27341_ (.A1(_16772_),
    .A2(_16771_),
    .ZN(_02177_));
 CLKBUF_X2 _27342_ (.A(_02177_),
    .Z(_02178_));
 NOR2_X2 _27343_ (.A1(_16774_),
    .A2(_16773_),
    .ZN(_02179_));
 AND2_X2 _27344_ (.A1(_02178_),
    .A2(_02179_),
    .ZN(_02180_));
 AOI221_X1 _27345_ (.A(_02172_),
    .B1(_02159_),
    .B2(_02173_),
    .C1(_02176_),
    .C2(_02180_),
    .ZN(_02181_));
 INV_X1 _27346_ (.A(_16769_),
    .ZN(_02182_));
 NOR2_X1 _27347_ (.A1(_02182_),
    .A2(_16770_),
    .ZN(_02183_));
 BUF_X2 _27348_ (.A(_02183_),
    .Z(_02184_));
 INV_X1 _27349_ (.A(_02184_),
    .ZN(_02185_));
 INV_X1 _27350_ (.A(_16768_),
    .ZN(_02186_));
 NOR2_X1 _27351_ (.A1(_02186_),
    .A2(_02158_),
    .ZN(_02187_));
 BUF_X2 _27352_ (.A(_02187_),
    .Z(_02188_));
 NOR2_X1 _27353_ (.A1(_02185_),
    .A2(_02188_),
    .ZN(_02189_));
 NAND2_X1 _27354_ (.A1(_02189_),
    .A2(_02151_),
    .ZN(_02190_));
 AND2_X2 _27355_ (.A1(_02168_),
    .A2(_02178_),
    .ZN(_02191_));
 BUF_X2 _27356_ (.A(_02191_),
    .Z(_02192_));
 AND2_X1 _27357_ (.A1(_02156_),
    .A2(_02166_),
    .ZN(_02193_));
 CLKBUF_X2 _27358_ (.A(_02193_),
    .Z(_02194_));
 AND2_X1 _27359_ (.A1(_02187_),
    .A2(_02142_),
    .ZN(_02195_));
 OR2_X1 _27360_ (.A1(_02194_),
    .A2(_02195_),
    .ZN(_02196_));
 NOR2_X1 _27361_ (.A1(_02163_),
    .A2(_16768_),
    .ZN(_02197_));
 CLKBUF_X2 _27362_ (.A(_02197_),
    .Z(_02198_));
 AND2_X1 _27363_ (.A1(_02198_),
    .A2(_02142_),
    .ZN(_02199_));
 BUF_X2 _27364_ (.A(_02199_),
    .Z(_02200_));
 OAI21_X1 _27365_ (.A(_02192_),
    .B1(_02196_),
    .B2(_02200_),
    .ZN(_02201_));
 AND4_X1 _27366_ (.A1(_02165_),
    .A2(_02181_),
    .A3(_02190_),
    .A4(_02201_),
    .ZN(_02202_));
 INV_X1 _27367_ (.A(_02193_),
    .ZN(_02203_));
 AND2_X1 _27368_ (.A1(_02157_),
    .A2(_02145_),
    .ZN(_02204_));
 INV_X1 _27369_ (.A(_02204_),
    .ZN(_02205_));
 NAND2_X1 _27370_ (.A1(_02203_),
    .A2(_02205_),
    .ZN(_02206_));
 NOR2_X1 _27371_ (.A1(_02169_),
    .A2(_16771_),
    .ZN(_02207_));
 AND2_X1 _27372_ (.A1(_02168_),
    .A2(_02207_),
    .ZN(_02208_));
 CLKBUF_X2 _27373_ (.A(_02208_),
    .Z(_02209_));
 AND2_X1 _27374_ (.A1(_02206_),
    .A2(_02209_),
    .ZN(_02210_));
 INV_X1 _27375_ (.A(_02210_),
    .ZN(_02211_));
 CLKBUF_X2 _27376_ (.A(_02173_),
    .Z(_02212_));
 INV_X1 _27377_ (.A(_02160_),
    .ZN(_02213_));
 NOR2_X1 _27378_ (.A1(_02213_),
    .A2(_02188_),
    .ZN(_02214_));
 BUF_X2 _27379_ (.A(_02209_),
    .Z(_02215_));
 AND2_X1 _27380_ (.A1(_02198_),
    .A2(_02157_),
    .ZN(_02216_));
 AOI22_X1 _27381_ (.A1(_02212_),
    .A2(_02214_),
    .B1(_02215_),
    .B2(_02216_),
    .ZN(_02217_));
 AND2_X1 _27382_ (.A1(_02211_),
    .A2(_02217_),
    .ZN(_02218_));
 AND2_X1 _27383_ (.A1(_02207_),
    .A2(_02148_),
    .ZN(_02219_));
 CLKBUF_X2 _27384_ (.A(_02219_),
    .Z(_02220_));
 BUF_X2 _27385_ (.A(_02167_),
    .Z(_02221_));
 AND2_X1 _27386_ (.A1(_02142_),
    .A2(_02186_),
    .ZN(_02222_));
 BUF_X2 _27387_ (.A(_02222_),
    .Z(_02223_));
 OAI21_X1 _27388_ (.A(_02220_),
    .B1(_02221_),
    .B2(_02223_),
    .ZN(_02224_));
 BUF_X2 _27389_ (.A(_02157_),
    .Z(_02225_));
 BUF_X2 _27390_ (.A(_02207_),
    .Z(_02226_));
 CLKBUF_X2 _27391_ (.A(_02148_),
    .Z(_02227_));
 NAND4_X1 _27392_ (.A1(_02198_),
    .A2(_02225_),
    .A3(_02226_),
    .A4(_02227_),
    .ZN(_02228_));
 NAND2_X1 _27393_ (.A1(_02224_),
    .A2(_02228_),
    .ZN(_02229_));
 INV_X1 _27394_ (.A(_02157_),
    .ZN(_02230_));
 NOR2_X1 _27395_ (.A1(_02230_),
    .A2(_02198_),
    .ZN(_02231_));
 AND2_X1 _27396_ (.A1(_16774_),
    .A2(_16773_),
    .ZN(_02232_));
 AND2_X1 _27397_ (.A1(_02226_),
    .A2(_02232_),
    .ZN(_02233_));
 BUF_X2 _27398_ (.A(_02233_),
    .Z(_02234_));
 BUF_X2 _27399_ (.A(_02234_),
    .Z(_02235_));
 AND2_X1 _27400_ (.A1(_02231_),
    .A2(_02235_),
    .ZN(_02236_));
 AND2_X1 _27401_ (.A1(_02148_),
    .A2(_02178_),
    .ZN(_02237_));
 CLKBUF_X2 _27402_ (.A(_02237_),
    .Z(_02238_));
 INV_X1 _27403_ (.A(_02188_),
    .ZN(_02239_));
 CLKBUF_X2 _27404_ (.A(_02184_),
    .Z(_02240_));
 AND3_X1 _27405_ (.A1(_02238_),
    .A2(_02239_),
    .A3(_02240_),
    .ZN(_02241_));
 NOR3_X1 _27406_ (.A1(_02229_),
    .A2(_02236_),
    .A3(_02241_),
    .ZN(_02242_));
 AND4_X1 _27407_ (.A1(_02154_),
    .A2(_02202_),
    .A3(_02218_),
    .A4(_02242_),
    .ZN(_02243_));
 AND2_X1 _27408_ (.A1(_02170_),
    .A2(_02232_),
    .ZN(_02244_));
 BUF_X2 _27409_ (.A(_02244_),
    .Z(_02245_));
 AND2_X2 _27410_ (.A1(_02197_),
    .A2(_02184_),
    .ZN(_02246_));
 AND2_X1 _27411_ (.A1(_02187_),
    .A2(_02161_),
    .ZN(_02247_));
 BUF_X2 _27412_ (.A(_02247_),
    .Z(_02248_));
 OAI21_X1 _27413_ (.A(_02245_),
    .B1(_02246_),
    .B2(_02248_),
    .ZN(_02249_));
 NAND2_X1 _27414_ (.A1(_02156_),
    .A2(_02186_),
    .ZN(_02250_));
 INV_X1 _27415_ (.A(_02250_),
    .ZN(_02251_));
 CLKBUF_X2 _27416_ (.A(_02251_),
    .Z(_02252_));
 NAND2_X1 _27417_ (.A1(_02244_),
    .A2(_02252_),
    .ZN(_02253_));
 AND2_X2 _27418_ (.A1(_02157_),
    .A2(_02187_),
    .ZN(_02254_));
 NAND2_X1 _27419_ (.A1(_02245_),
    .A2(_02254_),
    .ZN(_02255_));
 NAND2_X1 _27420_ (.A1(_02244_),
    .A2(_02194_),
    .ZN(_02256_));
 AND3_X1 _27421_ (.A1(_02253_),
    .A2(_02255_),
    .A3(_02256_),
    .ZN(_02257_));
 INV_X1 _27422_ (.A(_02166_),
    .ZN(_02258_));
 CLKBUF_X2 _27423_ (.A(_02258_),
    .Z(_02259_));
 CLKBUF_X2 _27424_ (.A(_02171_),
    .Z(_02260_));
 BUF_X2 _27425_ (.A(_02232_),
    .Z(_02261_));
 NAND4_X1 _27426_ (.A1(_02146_),
    .A2(_02259_),
    .A3(_02260_),
    .A4(_02261_),
    .ZN(_02262_));
 AND2_X1 _27427_ (.A1(_02232_),
    .A2(_02150_),
    .ZN(_02263_));
 CLKBUF_X2 _27428_ (.A(_02263_),
    .Z(_02264_));
 BUF_X2 _27429_ (.A(_02264_),
    .Z(_02265_));
 OAI21_X1 _27430_ (.A(_02265_),
    .B1(_02159_),
    .B2(_02223_),
    .ZN(_02266_));
 AND4_X1 _27431_ (.A1(_02249_),
    .A2(_02257_),
    .A3(_02262_),
    .A4(_02266_),
    .ZN(_02267_));
 AND2_X2 _27432_ (.A1(_02184_),
    .A2(_02186_),
    .ZN(_02268_));
 NAND2_X1 _27433_ (.A1(_02268_),
    .A2(_02234_),
    .ZN(_02269_));
 AND2_X1 _27434_ (.A1(_02177_),
    .A2(_02232_),
    .ZN(_02270_));
 CLKBUF_X2 _27435_ (.A(_16768_),
    .Z(_02271_));
 AND2_X1 _27436_ (.A1(_02161_),
    .A2(_02271_),
    .ZN(_02272_));
 AND2_X1 _27437_ (.A1(_02270_),
    .A2(_02272_),
    .ZN(_02273_));
 CLKBUF_X2 _27438_ (.A(_02270_),
    .Z(_02274_));
 CLKBUF_X2 _27439_ (.A(_02142_),
    .Z(_02275_));
 AND2_X1 _27440_ (.A1(_02275_),
    .A2(_02158_),
    .ZN(_02276_));
 AOI221_X4 _27441_ (.A(_02273_),
    .B1(_02225_),
    .B2(_02274_),
    .C1(_02234_),
    .C2(_02276_),
    .ZN(_02277_));
 NOR2_X2 _27442_ (.A1(_02213_),
    .A2(_02197_),
    .ZN(_02278_));
 NAND3_X1 _27443_ (.A1(_02235_),
    .A2(_02278_),
    .A3(_02239_),
    .ZN(_02279_));
 OAI21_X1 _27444_ (.A(_02155_),
    .B1(_02174_),
    .B2(_16769_),
    .ZN(_02280_));
 AND3_X1 _27445_ (.A1(_02150_),
    .A2(_02179_),
    .A3(_02155_),
    .ZN(_02281_));
 AND2_X1 _27446_ (.A1(_02280_),
    .A2(_02281_),
    .ZN(_02282_));
 INV_X1 _27447_ (.A(_02282_),
    .ZN(_02283_));
 BUF_X2 _27448_ (.A(_02168_),
    .Z(_02284_));
 BUF_X2 _27449_ (.A(_02158_),
    .Z(_02285_));
 NAND4_X1 _27450_ (.A1(_02284_),
    .A2(_02225_),
    .A3(_02285_),
    .A4(_02150_),
    .ZN(_02286_));
 AND2_X1 _27451_ (.A1(_02168_),
    .A2(_02150_),
    .ZN(_02287_));
 BUF_X2 _27452_ (.A(_02195_),
    .Z(_02288_));
 OAI21_X1 _27453_ (.A(_02287_),
    .B1(_02288_),
    .B2(_02223_),
    .ZN(_02289_));
 AND3_X1 _27454_ (.A1(_02283_),
    .A2(_02286_),
    .A3(_02289_),
    .ZN(_02290_));
 AND4_X1 _27455_ (.A1(_02269_),
    .A2(_02277_),
    .A3(_02279_),
    .A4(_02290_),
    .ZN(_02291_));
 AND2_X2 _27456_ (.A1(_02226_),
    .A2(_02179_),
    .ZN(_02292_));
 NAND2_X1 _27457_ (.A1(_02292_),
    .A2(_02247_),
    .ZN(_02293_));
 AND2_X1 _27458_ (.A1(_02161_),
    .A2(_02186_),
    .ZN(_02294_));
 NAND3_X1 _27459_ (.A1(_02294_),
    .A2(_02179_),
    .A3(_02226_),
    .ZN(_02295_));
 AND2_X1 _27460_ (.A1(_02293_),
    .A2(_02295_),
    .ZN(_02296_));
 AND2_X1 _27461_ (.A1(_02142_),
    .A2(_02145_),
    .ZN(_02297_));
 NOR2_X1 _27462_ (.A1(_02278_),
    .A2(_02297_),
    .ZN(_02298_));
 INV_X1 _27463_ (.A(_02237_),
    .ZN(_02299_));
 NOR2_X1 _27464_ (.A1(_02298_),
    .A2(_02299_),
    .ZN(_02300_));
 BUF_X2 _27465_ (.A(_02163_),
    .Z(_02301_));
 AND2_X1 _27466_ (.A1(_02263_),
    .A2(_02272_),
    .ZN(_02302_));
 AOI221_X4 _27467_ (.A(_02300_),
    .B1(_02301_),
    .B2(_02302_),
    .C1(_02288_),
    .C2(_02264_),
    .ZN(_02303_));
 AND2_X1 _27468_ (.A1(_02174_),
    .A2(_02157_),
    .ZN(_02304_));
 NAND2_X1 _27469_ (.A1(_02304_),
    .A2(_02292_),
    .ZN(_02305_));
 AND2_X1 _27470_ (.A1(_02197_),
    .A2(_02161_),
    .ZN(_02306_));
 AND2_X1 _27471_ (.A1(_02306_),
    .A2(_02270_),
    .ZN(_02307_));
 CLKBUF_X2 _27472_ (.A(_02274_),
    .Z(_02308_));
 AND2_X1 _27473_ (.A1(_02142_),
    .A2(_02163_),
    .ZN(_02309_));
 AND3_X1 _27474_ (.A1(_02308_),
    .A2(_02309_),
    .A3(_02271_),
    .ZN(_02310_));
 AND2_X2 _27475_ (.A1(_02183_),
    .A2(_02144_),
    .ZN(_02311_));
 AND2_X1 _27476_ (.A1(_02311_),
    .A2(_02274_),
    .ZN(_02312_));
 NOR3_X1 _27477_ (.A1(_02307_),
    .A2(_02310_),
    .A3(_02312_),
    .ZN(_02313_));
 AND4_X1 _27478_ (.A1(_02296_),
    .A2(_02303_),
    .A3(_02305_),
    .A4(_02313_),
    .ZN(_02314_));
 AND4_X1 _27479_ (.A1(_02243_),
    .A2(_02267_),
    .A3(_02291_),
    .A4(_02314_),
    .ZN(_02315_));
 AND2_X1 _27480_ (.A1(_02287_),
    .A2(_02311_),
    .ZN(_02316_));
 AND2_X1 _27481_ (.A1(_02166_),
    .A2(_02161_),
    .ZN(_02317_));
 CLKBUF_X2 _27482_ (.A(_02317_),
    .Z(_02318_));
 AND2_X1 _27483_ (.A1(_02215_),
    .A2(_02318_),
    .ZN(_02319_));
 AND2_X1 _27484_ (.A1(_02188_),
    .A2(_02184_),
    .ZN(_02320_));
 AND2_X1 _27485_ (.A1(_02209_),
    .A2(_02320_),
    .ZN(_02321_));
 AND2_X1 _27486_ (.A1(_02208_),
    .A2(_02306_),
    .ZN(_02322_));
 NOR4_X1 _27487_ (.A1(_02316_),
    .A2(_02319_),
    .A3(_02321_),
    .A4(_02322_),
    .ZN(_02323_));
 AND2_X1 _27488_ (.A1(_02170_),
    .A2(_02179_),
    .ZN(_02324_));
 BUF_X2 _27489_ (.A(_02324_),
    .Z(_02325_));
 CLKBUF_X2 _27490_ (.A(_02325_),
    .Z(_02326_));
 NOR3_X1 _27491_ (.A1(_02145_),
    .A2(_02182_),
    .A3(_16770_),
    .ZN(_02327_));
 AND2_X1 _27492_ (.A1(_02327_),
    .A2(_02258_),
    .ZN(_02328_));
 OAI21_X1 _27493_ (.A(_02326_),
    .B1(_02206_),
    .B2(_02328_),
    .ZN(_02329_));
 AND2_X1 _27494_ (.A1(_02171_),
    .A2(_02148_),
    .ZN(_02330_));
 AND4_X1 _27495_ (.A1(_02259_),
    .A2(_02330_),
    .A3(_02174_),
    .A4(_02162_),
    .ZN(_02331_));
 AND2_X1 _27496_ (.A1(_02142_),
    .A2(_02271_),
    .ZN(_02332_));
 BUF_X2 _27497_ (.A(_02332_),
    .Z(_02333_));
 BUF_X2 _27498_ (.A(_02330_),
    .Z(_02334_));
 AOI21_X1 _27499_ (.A(_02331_),
    .B1(_02333_),
    .B2(_02334_),
    .ZN(_02335_));
 AND2_X2 _27500_ (.A1(_02184_),
    .A2(_02158_),
    .ZN(_02336_));
 AND2_X2 _27501_ (.A1(_02161_),
    .A2(_02158_),
    .ZN(_02337_));
 OAI21_X1 _27502_ (.A(_02192_),
    .B1(_02336_),
    .B2(_02337_),
    .ZN(_02338_));
 BUF_X2 _27503_ (.A(_02292_),
    .Z(_02339_));
 OAI21_X1 _27504_ (.A(_02339_),
    .B1(_02328_),
    .B2(_02333_),
    .ZN(_02340_));
 AND4_X1 _27505_ (.A1(_02329_),
    .A2(_02335_),
    .A3(_02338_),
    .A4(_02340_),
    .ZN(_02341_));
 AND2_X1 _27506_ (.A1(_02209_),
    .A2(_02288_),
    .ZN(_02342_));
 INV_X1 _27507_ (.A(_02342_),
    .ZN(_02343_));
 AND2_X1 _27508_ (.A1(_02184_),
    .A2(_02166_),
    .ZN(_02344_));
 BUF_X2 _27509_ (.A(_02344_),
    .Z(_02345_));
 NAND2_X1 _27510_ (.A1(_02215_),
    .A2(_02345_),
    .ZN(_02346_));
 AND2_X2 _27511_ (.A1(_02145_),
    .A2(_02161_),
    .ZN(_02347_));
 AOI22_X1 _27512_ (.A1(_02192_),
    .A2(_02347_),
    .B1(_02220_),
    .B2(_02311_),
    .ZN(_02348_));
 NAND3_X1 _27513_ (.A1(_02343_),
    .A2(_02346_),
    .A3(_02348_),
    .ZN(_02349_));
 AND2_X1 _27514_ (.A1(_02149_),
    .A2(_02179_),
    .ZN(_02350_));
 BUF_X2 _27515_ (.A(_02350_),
    .Z(_02351_));
 BUF_X2 _27516_ (.A(_02225_),
    .Z(_02352_));
 BUF_X2 _27517_ (.A(_02184_),
    .Z(_02353_));
 OAI211_X1 _27518_ (.A(_02351_),
    .B(_02198_),
    .C1(_02352_),
    .C2(_02353_),
    .ZN(_02354_));
 INV_X1 _27519_ (.A(_02292_),
    .ZN(_02355_));
 BUF_X2 _27520_ (.A(_02297_),
    .Z(_02356_));
 INV_X1 _27521_ (.A(_02356_),
    .ZN(_02357_));
 BUF_X2 _27522_ (.A(_02180_),
    .Z(_02358_));
 INV_X1 _27523_ (.A(_02358_),
    .ZN(_02359_));
 OAI221_X1 _27524_ (.A(_02354_),
    .B1(_02355_),
    .B2(_02357_),
    .C1(_02205_),
    .C2(_02359_),
    .ZN(_02360_));
 BUF_X2 _27525_ (.A(_02272_),
    .Z(_02361_));
 AND2_X1 _27526_ (.A1(_02326_),
    .A2(_02361_),
    .ZN(_02362_));
 CLKBUF_X2 _27527_ (.A(_02320_),
    .Z(_02363_));
 INV_X1 _27528_ (.A(_02363_),
    .ZN(_02364_));
 INV_X1 _27529_ (.A(_02221_),
    .ZN(_02365_));
 AOI21_X1 _27530_ (.A(_02359_),
    .B1(_02364_),
    .B2(_02365_),
    .ZN(_02366_));
 NOR4_X1 _27531_ (.A1(_02349_),
    .A2(_02360_),
    .A3(_02362_),
    .A4(_02366_),
    .ZN(_02367_));
 AND2_X2 _27532_ (.A1(_02184_),
    .A2(_02271_),
    .ZN(_02368_));
 BUF_X2 _27533_ (.A(_02287_),
    .Z(_02369_));
 CLKBUF_X2 _27534_ (.A(_02294_),
    .Z(_02370_));
 AOI22_X1 _27535_ (.A1(_02212_),
    .A2(_02368_),
    .B1(_02369_),
    .B2(_02370_),
    .ZN(_02371_));
 NAND2_X1 _27536_ (.A1(_02209_),
    .A2(_02268_),
    .ZN(_02372_));
 INV_X1 _27537_ (.A(_02222_),
    .ZN(_02373_));
 OAI211_X1 _27538_ (.A(_02371_),
    .B(_02372_),
    .C1(_02373_),
    .C2(_02359_),
    .ZN(_02374_));
 BUF_X2 _27539_ (.A(_02186_),
    .Z(_02375_));
 INV_X1 _27540_ (.A(_02351_),
    .ZN(_02376_));
 AOI211_X1 _27541_ (.A(_02375_),
    .B(_02376_),
    .C1(_02213_),
    .C2(_02185_),
    .ZN(_02377_));
 AND2_X1 _27542_ (.A1(_02156_),
    .A2(_02271_),
    .ZN(_02378_));
 BUF_X2 _27543_ (.A(_02378_),
    .Z(_02379_));
 BUF_X2 _27544_ (.A(_02351_),
    .Z(_02380_));
 AND2_X1 _27545_ (.A1(_02379_),
    .A2(_02380_),
    .ZN(_02381_));
 AND3_X1 _27546_ (.A1(_02146_),
    .A2(_02259_),
    .A3(_02380_),
    .ZN(_02382_));
 NOR4_X1 _27547_ (.A1(_02374_),
    .A2(_02377_),
    .A3(_02381_),
    .A4(_02382_),
    .ZN(_02383_));
 AND4_X1 _27548_ (.A1(_02323_),
    .A2(_02341_),
    .A3(_02367_),
    .A4(_02383_),
    .ZN(_02384_));
 AND2_X2 _27549_ (.A1(_02315_),
    .A2(_02384_),
    .ZN(_02385_));
 INV_X1 _27550_ (.A(_16732_),
    .ZN(_02386_));
 AND2_X1 _27551_ (.A1(_02386_),
    .A2(_16731_),
    .ZN(_02387_));
 AND2_X1 _27552_ (.A1(_16734_),
    .A2(_16733_),
    .ZN(_02388_));
 CLKBUF_X2 _27553_ (.A(_02388_),
    .Z(_02389_));
 AND2_X1 _27554_ (.A1(_02387_),
    .A2(_02389_),
    .ZN(_02390_));
 CLKBUF_X2 _27555_ (.A(_02390_),
    .Z(_02391_));
 INV_X1 _27556_ (.A(_16729_),
    .ZN(_02392_));
 NOR2_X1 _27557_ (.A1(_02392_),
    .A2(_16730_),
    .ZN(_02393_));
 CLKBUF_X2 _27558_ (.A(_02393_),
    .Z(_02394_));
 INV_X1 _27559_ (.A(_16727_),
    .ZN(_02395_));
 NOR2_X1 _27560_ (.A1(_02395_),
    .A2(_16728_),
    .ZN(_02396_));
 CLKBUF_X2 _27561_ (.A(_02396_),
    .Z(_02397_));
 AND2_X2 _27562_ (.A1(_02394_),
    .A2(_02397_),
    .ZN(_02398_));
 INV_X1 _27563_ (.A(_16728_),
    .ZN(_02399_));
 NOR2_X1 _27564_ (.A1(_02399_),
    .A2(_16727_),
    .ZN(_02400_));
 CLKBUF_X2 _27565_ (.A(_02400_),
    .Z(_02401_));
 NOR2_X1 _27566_ (.A1(_16729_),
    .A2(_16730_),
    .ZN(_02402_));
 CLKBUF_X2 _27567_ (.A(_02402_),
    .Z(_02403_));
 AND2_X2 _27568_ (.A1(_02401_),
    .A2(_02403_),
    .ZN(_02404_));
 NOR2_X1 _27569_ (.A1(_02398_),
    .A2(_02404_),
    .ZN(_02405_));
 INV_X1 _27570_ (.A(_02405_),
    .ZN(_02406_));
 AND2_X2 _27571_ (.A1(_16729_),
    .A2(_16730_),
    .ZN(_02407_));
 AND2_X2 _27572_ (.A1(_02397_),
    .A2(_02407_),
    .ZN(_02408_));
 INV_X1 _27573_ (.A(_02408_),
    .ZN(_02409_));
 AND2_X2 _27574_ (.A1(_02401_),
    .A2(_02407_),
    .ZN(_02410_));
 INV_X1 _27575_ (.A(_02410_),
    .ZN(_02411_));
 INV_X1 _27576_ (.A(_16730_),
    .ZN(_02412_));
 NOR2_X2 _27577_ (.A1(_02412_),
    .A2(_16729_),
    .ZN(_02413_));
 INV_X1 _27578_ (.A(_02413_),
    .ZN(_02414_));
 NAND3_X1 _27579_ (.A1(_02409_),
    .A2(_02411_),
    .A3(_02414_),
    .ZN(_02415_));
 OAI21_X1 _27580_ (.A(_02391_),
    .B1(_02406_),
    .B2(_02415_),
    .ZN(_02416_));
 NOR2_X2 _27581_ (.A1(_16732_),
    .A2(_16731_),
    .ZN(_02417_));
 AND2_X1 _27582_ (.A1(_02388_),
    .A2(_02417_),
    .ZN(_02418_));
 INV_X2 _27583_ (.A(_02418_),
    .ZN(_02419_));
 AND2_X1 _27584_ (.A1(_02397_),
    .A2(_02413_),
    .ZN(_02420_));
 INV_X1 _27585_ (.A(_02420_),
    .ZN(_02421_));
 AND2_X1 _27586_ (.A1(_16728_),
    .A2(_16727_),
    .ZN(_02422_));
 CLKBUF_X2 _27587_ (.A(_02422_),
    .Z(_02423_));
 AND2_X1 _27588_ (.A1(_02413_),
    .A2(_02423_),
    .ZN(_02424_));
 INV_X1 _27589_ (.A(_02424_),
    .ZN(_02425_));
 AOI21_X1 _27590_ (.A(_02419_),
    .B1(_02421_),
    .B2(_02425_),
    .ZN(_02426_));
 INV_X1 _27591_ (.A(_02407_),
    .ZN(_02427_));
 CLKBUF_X2 _27592_ (.A(_16728_),
    .Z(_02428_));
 CLKBUF_X2 _27593_ (.A(_16727_),
    .Z(_02429_));
 BUF_X2 _27594_ (.A(_02429_),
    .Z(_02430_));
 AOI211_X1 _27595_ (.A(_02427_),
    .B(_02419_),
    .C1(_02428_),
    .C2(_02430_),
    .ZN(_02431_));
 BUF_X2 _27596_ (.A(_02418_),
    .Z(_02432_));
 AOI211_X1 _27597_ (.A(_02426_),
    .B(_02431_),
    .C1(_02404_),
    .C2(_02432_),
    .ZN(_02433_));
 CLKBUF_X2 _27598_ (.A(_02413_),
    .Z(_02434_));
 BUF_X2 _27599_ (.A(_02434_),
    .Z(_02435_));
 NOR2_X2 _27600_ (.A1(_02386_),
    .A2(_16731_),
    .ZN(_02436_));
 BUF_X2 _27601_ (.A(_02436_),
    .Z(_02437_));
 CLKBUF_X2 _27602_ (.A(_02389_),
    .Z(_02438_));
 NAND4_X1 _27603_ (.A1(_02435_),
    .A2(_02437_),
    .A3(_02428_),
    .A4(_02438_),
    .ZN(_02439_));
 AND2_X1 _27604_ (.A1(_02436_),
    .A2(_02388_),
    .ZN(_02440_));
 CLKBUF_X2 _27605_ (.A(_02440_),
    .Z(_02441_));
 BUF_X2 _27606_ (.A(_02441_),
    .Z(_02442_));
 AND2_X1 _27607_ (.A1(_02422_),
    .A2(_02402_),
    .ZN(_02443_));
 INV_X1 _27608_ (.A(_02443_),
    .ZN(_02444_));
 NOR2_X1 _27609_ (.A1(_16728_),
    .A2(_16727_),
    .ZN(_02445_));
 AND2_X1 _27610_ (.A1(_02402_),
    .A2(_02445_),
    .ZN(_02446_));
 INV_X1 _27611_ (.A(_02446_),
    .ZN(_02447_));
 NAND2_X1 _27612_ (.A1(_02444_),
    .A2(_02447_),
    .ZN(_02448_));
 AND2_X1 _27613_ (.A1(_02393_),
    .A2(_02399_),
    .ZN(_02449_));
 BUF_X2 _27614_ (.A(_02449_),
    .Z(_02450_));
 OAI21_X1 _27615_ (.A(_02442_),
    .B1(_02448_),
    .B2(_02450_),
    .ZN(_02451_));
 BUF_X2 _27616_ (.A(_02445_),
    .Z(_02452_));
 NAND4_X1 _27617_ (.A1(_02435_),
    .A2(_02437_),
    .A3(_02438_),
    .A4(_02452_),
    .ZN(_02453_));
 CLKBUF_X2 _27618_ (.A(_02407_),
    .Z(_02454_));
 AND2_X1 _27619_ (.A1(_02454_),
    .A2(_16727_),
    .ZN(_02455_));
 NAND3_X1 _27620_ (.A1(_02455_),
    .A2(_02438_),
    .A3(_02437_),
    .ZN(_02456_));
 AND4_X1 _27621_ (.A1(_02439_),
    .A2(_02451_),
    .A3(_02453_),
    .A4(_02456_),
    .ZN(_02457_));
 AND2_X1 _27622_ (.A1(_02393_),
    .A2(_02445_),
    .ZN(_02458_));
 AND2_X2 _27623_ (.A1(_16732_),
    .A2(_16731_),
    .ZN(_02459_));
 AND2_X1 _27624_ (.A1(_02388_),
    .A2(_02459_),
    .ZN(_02460_));
 BUF_X2 _27625_ (.A(_02460_),
    .Z(_02461_));
 BUF_X2 _27626_ (.A(_02461_),
    .Z(_02462_));
 NAND2_X1 _27627_ (.A1(_02458_),
    .A2(_02462_),
    .ZN(_02463_));
 NOR2_X1 _27628_ (.A1(_02412_),
    .A2(_16728_),
    .ZN(_02464_));
 AND2_X1 _27629_ (.A1(_02464_),
    .A2(_02392_),
    .ZN(_02465_));
 BUF_X2 _27630_ (.A(_02465_),
    .Z(_02466_));
 AND2_X2 _27631_ (.A1(_02413_),
    .A2(_16728_),
    .ZN(_02467_));
 BUF_X2 _27632_ (.A(_02467_),
    .Z(_02468_));
 OAI21_X1 _27633_ (.A(_02462_),
    .B1(_02466_),
    .B2(_02468_),
    .ZN(_02469_));
 CLKBUF_X2 _27634_ (.A(_02403_),
    .Z(_02470_));
 OAI211_X1 _27635_ (.A(_02462_),
    .B(_02470_),
    .C1(_02428_),
    .C2(_02430_),
    .ZN(_02471_));
 CLKBUF_X2 _27636_ (.A(_02401_),
    .Z(_02472_));
 NAND3_X1 _27637_ (.A1(_02461_),
    .A2(_02472_),
    .A3(_02454_),
    .ZN(_02473_));
 AND4_X1 _27638_ (.A1(_02463_),
    .A2(_02469_),
    .A3(_02471_),
    .A4(_02473_),
    .ZN(_02474_));
 AND4_X1 _27639_ (.A1(_02416_),
    .A2(_02433_),
    .A3(_02457_),
    .A4(_02474_),
    .ZN(_02475_));
 AND2_X2 _27640_ (.A1(_02422_),
    .A2(_02407_),
    .ZN(_02476_));
 NOR2_X1 _27641_ (.A1(_16734_),
    .A2(_16733_),
    .ZN(_02477_));
 AND2_X1 _27642_ (.A1(_02459_),
    .A2(_02477_),
    .ZN(_02478_));
 CLKBUF_X2 _27643_ (.A(_02478_),
    .Z(_02479_));
 AND2_X1 _27644_ (.A1(_02476_),
    .A2(_02479_),
    .ZN(_02480_));
 AND2_X1 _27645_ (.A1(_02407_),
    .A2(_02399_),
    .ZN(_02481_));
 AND2_X1 _27646_ (.A1(_02481_),
    .A2(_02478_),
    .ZN(_02482_));
 AND2_X1 _27647_ (.A1(_02413_),
    .A2(_02452_),
    .ZN(_02483_));
 AOI211_X1 _27648_ (.A(_02480_),
    .B(_02482_),
    .C1(_02479_),
    .C2(_02483_),
    .ZN(_02484_));
 INV_X1 _27649_ (.A(_02403_),
    .ZN(_02485_));
 NOR2_X1 _27650_ (.A1(_02485_),
    .A2(_02452_),
    .ZN(_02486_));
 NAND2_X1 _27651_ (.A1(_02486_),
    .A2(_02478_),
    .ZN(_02487_));
 INV_X1 _27652_ (.A(_02478_),
    .ZN(_02488_));
 AND2_X1 _27653_ (.A1(_02401_),
    .A2(_02393_),
    .ZN(_02489_));
 INV_X1 _27654_ (.A(_02489_),
    .ZN(_02490_));
 OAI211_X1 _27655_ (.A(_02484_),
    .B(_02487_),
    .C1(_02488_),
    .C2(_02490_),
    .ZN(_02491_));
 AND2_X1 _27656_ (.A1(_02417_),
    .A2(_02477_),
    .ZN(_02492_));
 CLKBUF_X2 _27657_ (.A(_02492_),
    .Z(_02493_));
 AND2_X1 _27658_ (.A1(_02402_),
    .A2(_16728_),
    .ZN(_02494_));
 BUF_X2 _27659_ (.A(_02494_),
    .Z(_02495_));
 AND2_X1 _27660_ (.A1(_02493_),
    .A2(_02495_),
    .ZN(_02496_));
 AND3_X1 _27661_ (.A1(_02493_),
    .A2(_02394_),
    .A3(_02397_),
    .ZN(_02497_));
 BUF_X2 _27662_ (.A(_02493_),
    .Z(_02498_));
 AND2_X1 _27663_ (.A1(_02393_),
    .A2(_16728_),
    .ZN(_02499_));
 BUF_X2 _27664_ (.A(_02499_),
    .Z(_02500_));
 AOI211_X1 _27665_ (.A(_02496_),
    .B(_02497_),
    .C1(_02498_),
    .C2(_02500_),
    .ZN(_02501_));
 OR2_X1 _27666_ (.A1(_02424_),
    .A2(_02483_),
    .ZN(_02502_));
 AND2_X1 _27667_ (.A1(_02387_),
    .A2(_02477_),
    .ZN(_02503_));
 BUF_X2 _27668_ (.A(_02503_),
    .Z(_02504_));
 NAND2_X1 _27669_ (.A1(_02502_),
    .A2(_02504_),
    .ZN(_02505_));
 INV_X1 _27670_ (.A(_02445_),
    .ZN(_02506_));
 AND2_X1 _27671_ (.A1(_02506_),
    .A2(_02394_),
    .ZN(_02507_));
 INV_X1 _27672_ (.A(_02423_),
    .ZN(_02508_));
 AND2_X1 _27673_ (.A1(_02507_),
    .A2(_02508_),
    .ZN(_02509_));
 OAI21_X1 _27674_ (.A(_02504_),
    .B1(_02509_),
    .B2(_02495_),
    .ZN(_02510_));
 NOR2_X1 _27675_ (.A1(_02427_),
    .A2(_02423_),
    .ZN(_02511_));
 OAI221_X1 _27676_ (.A(_02498_),
    .B1(_02428_),
    .B2(_02430_),
    .C1(_02511_),
    .C2(_02435_),
    .ZN(_02512_));
 NAND4_X1 _27677_ (.A1(_02501_),
    .A2(_02505_),
    .A3(_02510_),
    .A4(_02512_),
    .ZN(_02513_));
 AND2_X1 _27678_ (.A1(_02436_),
    .A2(_02477_),
    .ZN(_02514_));
 BUF_X2 _27679_ (.A(_02514_),
    .Z(_02515_));
 INV_X1 _27680_ (.A(_02515_),
    .ZN(_02516_));
 INV_X1 _27681_ (.A(_02507_),
    .ZN(_02517_));
 AOI211_X1 _27682_ (.A(_02423_),
    .B(_02516_),
    .C1(_02485_),
    .C2(_02517_),
    .ZN(_02518_));
 AND2_X1 _27683_ (.A1(_02506_),
    .A2(_02413_),
    .ZN(_02519_));
 AND2_X1 _27684_ (.A1(_02519_),
    .A2(_02514_),
    .ZN(_02520_));
 INV_X1 _27685_ (.A(_02520_),
    .ZN(_02521_));
 AND2_X1 _27686_ (.A1(_02407_),
    .A2(_02428_),
    .ZN(_02522_));
 BUF_X2 _27687_ (.A(_02522_),
    .Z(_02523_));
 CLKBUF_X2 _27688_ (.A(_02477_),
    .Z(_02524_));
 NAND3_X1 _27689_ (.A1(_02523_),
    .A2(_02437_),
    .A3(_02524_),
    .ZN(_02525_));
 AND2_X1 _27690_ (.A1(_02407_),
    .A2(_02445_),
    .ZN(_02526_));
 CLKBUF_X2 _27691_ (.A(_02526_),
    .Z(_02527_));
 INV_X1 _27692_ (.A(_02527_),
    .ZN(_02528_));
 OAI211_X1 _27693_ (.A(_02521_),
    .B(_02525_),
    .C1(_02528_),
    .C2(_02516_),
    .ZN(_02529_));
 NOR4_X1 _27694_ (.A1(_02491_),
    .A2(_02513_),
    .A3(_02518_),
    .A4(_02529_),
    .ZN(_02530_));
 INV_X1 _27695_ (.A(_16734_),
    .ZN(_02531_));
 NOR2_X2 _27696_ (.A1(_02531_),
    .A2(_16733_),
    .ZN(_02532_));
 AND2_X1 _27697_ (.A1(_02387_),
    .A2(_02532_),
    .ZN(_02533_));
 CLKBUF_X2 _27698_ (.A(_02533_),
    .Z(_02534_));
 AND3_X1 _27699_ (.A1(_02534_),
    .A2(_02508_),
    .A3(_02486_),
    .ZN(_02535_));
 AOI21_X1 _27700_ (.A(_02535_),
    .B1(_02534_),
    .B2(_02523_),
    .ZN(_02536_));
 AND2_X1 _27701_ (.A1(_02436_),
    .A2(_02532_),
    .ZN(_02537_));
 AND2_X1 _27702_ (.A1(_02537_),
    .A2(_02476_),
    .ZN(_02538_));
 INV_X1 _27703_ (.A(_02538_),
    .ZN(_02539_));
 BUF_X2 _27704_ (.A(_02537_),
    .Z(_02540_));
 BUF_X2 _27705_ (.A(_02481_),
    .Z(_02541_));
 OAI21_X1 _27706_ (.A(_02540_),
    .B1(_02420_),
    .B2(_02541_),
    .ZN(_02542_));
 INV_X1 _27707_ (.A(_02540_),
    .ZN(_02543_));
 INV_X1 _27708_ (.A(_02458_),
    .ZN(_02544_));
 OAI211_X1 _27709_ (.A(_02539_),
    .B(_02542_),
    .C1(_02543_),
    .C2(_02544_),
    .ZN(_02545_));
 INV_X1 _27710_ (.A(_02393_),
    .ZN(_02546_));
 NOR2_X1 _27711_ (.A1(_02546_),
    .A2(_02401_),
    .ZN(_02547_));
 AND2_X1 _27712_ (.A1(_02532_),
    .A2(_02459_),
    .ZN(_02548_));
 BUF_X2 _27713_ (.A(_02548_),
    .Z(_02549_));
 AND2_X1 _27714_ (.A1(_02547_),
    .A2(_02549_),
    .ZN(_02550_));
 NOR2_X1 _27715_ (.A1(_02485_),
    .A2(_02397_),
    .ZN(_02551_));
 AND2_X1 _27716_ (.A1(_02549_),
    .A2(_02551_),
    .ZN(_02552_));
 CLKBUF_X2 _27717_ (.A(_02532_),
    .Z(_02553_));
 CLKBUF_X2 _27718_ (.A(_02459_),
    .Z(_02554_));
 AND3_X1 _27719_ (.A1(_02527_),
    .A2(_02553_),
    .A3(_02554_),
    .ZN(_02555_));
 NOR4_X1 _27720_ (.A1(_02545_),
    .A2(_02550_),
    .A3(_02552_),
    .A4(_02555_),
    .ZN(_02556_));
 CLKBUF_X2 _27721_ (.A(_02395_),
    .Z(_02557_));
 CLKBUF_X2 _27722_ (.A(_02417_),
    .Z(_02558_));
 AND4_X1 _27723_ (.A1(_02557_),
    .A2(_02553_),
    .A3(_02470_),
    .A4(_02558_),
    .ZN(_02559_));
 AND2_X2 _27724_ (.A1(_02532_),
    .A2(_02417_),
    .ZN(_02560_));
 BUF_X2 _27725_ (.A(_02560_),
    .Z(_02561_));
 AOI21_X1 _27726_ (.A(_02559_),
    .B1(_02561_),
    .B2(_02547_),
    .ZN(_02562_));
 NOR2_X1 _27727_ (.A1(_02427_),
    .A2(_02452_),
    .ZN(_02563_));
 AND2_X1 _27728_ (.A1(_02434_),
    .A2(_02429_),
    .ZN(_02564_));
 OAI21_X1 _27729_ (.A(_02561_),
    .B1(_02563_),
    .B2(_02564_),
    .ZN(_02565_));
 AND4_X1 _27730_ (.A1(_02536_),
    .A2(_02556_),
    .A3(_02562_),
    .A4(_02565_),
    .ZN(_02566_));
 AND2_X1 _27731_ (.A1(_02531_),
    .A2(_16733_),
    .ZN(_02567_));
 AND2_X1 _27732_ (.A1(_02567_),
    .A2(_02417_),
    .ZN(_02568_));
 INV_X1 _27733_ (.A(_02568_),
    .ZN(_02569_));
 AND2_X1 _27734_ (.A1(_02403_),
    .A2(_02399_),
    .ZN(_02570_));
 BUF_X2 _27735_ (.A(_02570_),
    .Z(_02571_));
 INV_X1 _27736_ (.A(_02571_),
    .ZN(_02572_));
 AOI21_X1 _27737_ (.A(_02569_),
    .B1(_02544_),
    .B2(_02572_),
    .ZN(_02573_));
 AND2_X1 _27738_ (.A1(_02567_),
    .A2(_02387_),
    .ZN(_02574_));
 BUF_X2 _27739_ (.A(_02574_),
    .Z(_02575_));
 NAND2_X1 _27740_ (.A1(_02575_),
    .A2(_02500_),
    .ZN(_02576_));
 NAND2_X1 _27741_ (.A1(_02575_),
    .A2(_02571_),
    .ZN(_02577_));
 BUF_X2 _27742_ (.A(_02443_),
    .Z(_02578_));
 NAND2_X1 _27743_ (.A1(_02575_),
    .A2(_02578_),
    .ZN(_02579_));
 NAND3_X1 _27744_ (.A1(_02576_),
    .A2(_02577_),
    .A3(_02579_),
    .ZN(_02580_));
 BUF_X2 _27745_ (.A(_02568_),
    .Z(_02581_));
 OAI21_X1 _27746_ (.A(_02581_),
    .B1(_02410_),
    .B2(_02541_),
    .ZN(_02582_));
 CLKBUF_X2 _27747_ (.A(_02567_),
    .Z(_02583_));
 NAND4_X1 _27748_ (.A1(_02583_),
    .A2(_02429_),
    .A3(_02434_),
    .A4(_02558_),
    .ZN(_02584_));
 NAND2_X1 _27749_ (.A1(_02582_),
    .A2(_02584_),
    .ZN(_02585_));
 CLKBUF_X2 _27750_ (.A(_02387_),
    .Z(_02586_));
 NAND4_X1 _27751_ (.A1(_02583_),
    .A2(_02586_),
    .A3(_02434_),
    .A4(_02429_),
    .ZN(_02587_));
 INV_X1 _27752_ (.A(_02575_),
    .ZN(_02588_));
 INV_X1 _27753_ (.A(_02476_),
    .ZN(_02589_));
 OAI21_X1 _27754_ (.A(_02587_),
    .B1(_02588_),
    .B2(_02589_),
    .ZN(_02590_));
 OR4_X1 _27755_ (.A1(_02573_),
    .A2(_02580_),
    .A3(_02585_),
    .A4(_02590_),
    .ZN(_02591_));
 AND2_X1 _27756_ (.A1(_02567_),
    .A2(_02459_),
    .ZN(_02592_));
 BUF_X2 _27757_ (.A(_02592_),
    .Z(_02593_));
 NAND3_X1 _27758_ (.A1(_02593_),
    .A2(_02508_),
    .A3(_02563_),
    .ZN(_02594_));
 BUF_X2 _27759_ (.A(_02424_),
    .Z(_02595_));
 BUF_X2 _27760_ (.A(_02583_),
    .Z(_02596_));
 NAND3_X1 _27761_ (.A1(_02595_),
    .A2(_02596_),
    .A3(_02554_),
    .ZN(_02597_));
 NAND2_X1 _27762_ (.A1(_02594_),
    .A2(_02597_),
    .ZN(_02598_));
 AND2_X2 _27763_ (.A1(_02567_),
    .A2(_02436_),
    .ZN(_02599_));
 BUF_X2 _27764_ (.A(_02599_),
    .Z(_02600_));
 OAI21_X1 _27765_ (.A(_02600_),
    .B1(_02500_),
    .B2(_02450_),
    .ZN(_02601_));
 AND2_X2 _27766_ (.A1(_02396_),
    .A2(_02403_),
    .ZN(_02602_));
 OAI21_X1 _27767_ (.A(_02600_),
    .B1(_02602_),
    .B2(_02578_),
    .ZN(_02603_));
 NAND2_X1 _27768_ (.A1(_02599_),
    .A2(_02410_),
    .ZN(_02604_));
 NOR2_X1 _27769_ (.A1(_02414_),
    .A2(_02401_),
    .ZN(_02605_));
 NAND2_X1 _27770_ (.A1(_02605_),
    .A2(_02599_),
    .ZN(_02606_));
 NAND4_X1 _27771_ (.A1(_02601_),
    .A2(_02603_),
    .A3(_02604_),
    .A4(_02606_),
    .ZN(_02607_));
 NAND2_X1 _27772_ (.A1(_02592_),
    .A2(_02443_),
    .ZN(_02608_));
 NOR2_X1 _27773_ (.A1(_02395_),
    .A2(_16730_),
    .ZN(_02609_));
 AND2_X1 _27774_ (.A1(_02609_),
    .A2(_16729_),
    .ZN(_02610_));
 NAND3_X1 _27775_ (.A1(_02610_),
    .A2(_02596_),
    .A3(_02554_),
    .ZN(_02611_));
 INV_X1 _27776_ (.A(_02593_),
    .ZN(_02612_));
 OAI211_X1 _27777_ (.A(_02608_),
    .B(_02611_),
    .C1(_02612_),
    .C2(_02572_),
    .ZN(_02613_));
 NOR4_X1 _27778_ (.A1(_02591_),
    .A2(_02598_),
    .A3(_02607_),
    .A4(_02613_),
    .ZN(_02614_));
 NAND4_X1 _27779_ (.A1(_02475_),
    .A2(_02530_),
    .A3(_02566_),
    .A4(_02614_),
    .ZN(_02615_));
 AND2_X1 _27780_ (.A1(_02498_),
    .A2(_02446_),
    .ZN(_02616_));
 OR2_X2 _27781_ (.A1(_02615_),
    .A2(_02616_),
    .ZN(_02617_));
 XNOR2_X1 _27782_ (.A(_02385_),
    .B(_02617_),
    .ZN(_02618_));
 XNOR2_X1 _27783_ (.A(_02141_),
    .B(_02618_),
    .ZN(_02619_));
 INV_X1 _27784_ (.A(_16782_),
    .ZN(_02620_));
 AND2_X1 _27785_ (.A1(_02620_),
    .A2(_16781_),
    .ZN(_02621_));
 CLKBUF_X2 _27786_ (.A(_02621_),
    .Z(_02622_));
 AND2_X1 _27787_ (.A1(_16780_),
    .A2(_16779_),
    .ZN(_02623_));
 AND2_X1 _27788_ (.A1(_02622_),
    .A2(_02623_),
    .ZN(_02624_));
 INV_X1 _27789_ (.A(_16776_),
    .ZN(_02625_));
 BUF_X2 _27790_ (.A(_16775_),
    .Z(_02626_));
 NOR2_X2 _27791_ (.A1(_02625_),
    .A2(_02626_),
    .ZN(_02627_));
 INV_X1 _27792_ (.A(_16778_),
    .ZN(_02628_));
 NOR2_X2 _27793_ (.A1(_02628_),
    .A2(_16777_),
    .ZN(_02629_));
 AND2_X1 _27794_ (.A1(_02627_),
    .A2(_02629_),
    .ZN(_02630_));
 AND2_X1 _27795_ (.A1(_02624_),
    .A2(_02630_),
    .ZN(_02631_));
 AND2_X1 _27796_ (.A1(_02629_),
    .A2(_02625_),
    .ZN(_02632_));
 AND2_X1 _27797_ (.A1(_02624_),
    .A2(_02632_),
    .ZN(_02633_));
 NOR2_X1 _27798_ (.A1(_02631_),
    .A2(_02633_),
    .ZN(_02634_));
 BUF_X2 _27799_ (.A(_02624_),
    .Z(_02635_));
 INV_X1 _27800_ (.A(_16775_),
    .ZN(_02636_));
 NOR2_X1 _27801_ (.A1(_02636_),
    .A2(_16776_),
    .ZN(_02637_));
 CLKBUF_X2 _27802_ (.A(_02637_),
    .Z(_02638_));
 AND2_X1 _27803_ (.A1(_16777_),
    .A2(_16778_),
    .ZN(_02639_));
 AND2_X1 _27804_ (.A1(_02638_),
    .A2(_02639_),
    .ZN(_02640_));
 BUF_X2 _27805_ (.A(_02640_),
    .Z(_02641_));
 BUF_X2 _27806_ (.A(_16776_),
    .Z(_02642_));
 AND2_X1 _27807_ (.A1(_02639_),
    .A2(_02642_),
    .ZN(_02643_));
 OAI21_X1 _27808_ (.A(_02635_),
    .B1(_02641_),
    .B2(_02643_),
    .ZN(_02644_));
 AND2_X1 _27809_ (.A1(_02634_),
    .A2(_02644_),
    .ZN(_02645_));
 NOR2_X1 _27810_ (.A1(_16777_),
    .A2(_16778_),
    .ZN(_02646_));
 AND2_X1 _27811_ (.A1(_02646_),
    .A2(_02626_),
    .ZN(_02647_));
 AND2_X1 _27812_ (.A1(_02624_),
    .A2(_02647_),
    .ZN(_02648_));
 INV_X1 _27813_ (.A(_02648_),
    .ZN(_02649_));
 INV_X1 _27814_ (.A(_16777_),
    .ZN(_02650_));
 NOR2_X1 _27815_ (.A1(_02650_),
    .A2(_16778_),
    .ZN(_02651_));
 AND2_X1 _27816_ (.A1(_16775_),
    .A2(_16776_),
    .ZN(_02652_));
 AND2_X1 _27817_ (.A1(_02651_),
    .A2(_02652_),
    .ZN(_02653_));
 BUF_X2 _27818_ (.A(_02653_),
    .Z(_02654_));
 NAND2_X1 _27819_ (.A1(_02624_),
    .A2(_02654_),
    .ZN(_02655_));
 CLKBUF_X2 _27820_ (.A(_02651_),
    .Z(_02656_));
 BUF_X2 _27821_ (.A(_02625_),
    .Z(_02657_));
 AND2_X2 _27822_ (.A1(_02656_),
    .A2(_02657_),
    .ZN(_02658_));
 NAND2_X1 _27823_ (.A1(_02624_),
    .A2(_02658_),
    .ZN(_02659_));
 AND3_X1 _27824_ (.A1(_02649_),
    .A2(_02655_),
    .A3(_02659_),
    .ZN(_02660_));
 INV_X1 _27825_ (.A(_16780_),
    .ZN(_02661_));
 NOR2_X2 _27826_ (.A1(_02661_),
    .A2(_16779_),
    .ZN(_02662_));
 AND2_X1 _27827_ (.A1(_02621_),
    .A2(_02662_),
    .ZN(_02663_));
 CLKBUF_X2 _27828_ (.A(_02663_),
    .Z(_02664_));
 BUF_X2 _27829_ (.A(_02664_),
    .Z(_02665_));
 CLKBUF_X2 _27830_ (.A(_02646_),
    .Z(_02666_));
 BUF_X2 _27831_ (.A(_02666_),
    .Z(_02667_));
 OAI21_X1 _27832_ (.A(_02665_),
    .B1(_02654_),
    .B2(_02667_),
    .ZN(_02668_));
 AND2_X1 _27833_ (.A1(_02637_),
    .A2(_02629_),
    .ZN(_02669_));
 BUF_X2 _27834_ (.A(_02669_),
    .Z(_02670_));
 BUF_X2 _27835_ (.A(_02643_),
    .Z(_02671_));
 OAI21_X1 _27836_ (.A(_02665_),
    .B1(_02670_),
    .B2(_02671_),
    .ZN(_02672_));
 AND4_X1 _27837_ (.A1(_02645_),
    .A2(_02660_),
    .A3(_02668_),
    .A4(_02672_),
    .ZN(_02673_));
 CLKBUF_X2 _27838_ (.A(_02639_),
    .Z(_02674_));
 AND2_X2 _27839_ (.A1(_02674_),
    .A2(_02657_),
    .ZN(_02675_));
 NOR2_X2 _27840_ (.A1(_16780_),
    .A2(_16779_),
    .ZN(_02676_));
 NOR2_X1 _27841_ (.A1(_16782_),
    .A2(_16781_),
    .ZN(_02677_));
 CLKBUF_X2 _27842_ (.A(_02677_),
    .Z(_02678_));
 AND2_X1 _27843_ (.A1(_02676_),
    .A2(_02678_),
    .ZN(_02679_));
 BUF_X2 _27844_ (.A(_02679_),
    .Z(_02680_));
 NAND2_X1 _27845_ (.A1(_02675_),
    .A2(_02680_),
    .ZN(_02681_));
 AND2_X1 _27846_ (.A1(_02627_),
    .A2(_02674_),
    .ZN(_02682_));
 NAND2_X1 _27847_ (.A1(_02682_),
    .A2(_02680_),
    .ZN(_02683_));
 NOR2_X2 _27848_ (.A1(_02626_),
    .A2(_16776_),
    .ZN(_02684_));
 AND2_X1 _27849_ (.A1(_02656_),
    .A2(_02684_),
    .ZN(_02685_));
 BUF_X2 _27850_ (.A(_02685_),
    .Z(_02686_));
 INV_X1 _27851_ (.A(_02686_),
    .ZN(_02687_));
 INV_X1 _27852_ (.A(_02654_),
    .ZN(_02688_));
 NAND2_X1 _27853_ (.A1(_02687_),
    .A2(_02688_),
    .ZN(_02689_));
 INV_X1 _27854_ (.A(_02689_),
    .ZN(_02690_));
 INV_X1 _27855_ (.A(_02680_),
    .ZN(_02691_));
 OAI211_X1 _27856_ (.A(_02681_),
    .B(_02683_),
    .C1(_02690_),
    .C2(_02691_),
    .ZN(_02692_));
 INV_X1 _27857_ (.A(_16779_),
    .ZN(_02693_));
 NOR2_X2 _27858_ (.A1(_02693_),
    .A2(_16780_),
    .ZN(_02694_));
 AND2_X2 _27859_ (.A1(_02694_),
    .A2(_02678_),
    .ZN(_02695_));
 AND2_X2 _27860_ (.A1(_02646_),
    .A2(_02625_),
    .ZN(_02696_));
 NAND2_X1 _27861_ (.A1(_02695_),
    .A2(_02696_),
    .ZN(_02697_));
 AND2_X2 _27862_ (.A1(_02627_),
    .A2(_02646_),
    .ZN(_02698_));
 NAND2_X1 _27863_ (.A1(_02698_),
    .A2(_02695_),
    .ZN(_02699_));
 INV_X1 _27864_ (.A(_02695_),
    .ZN(_02700_));
 OAI211_X1 _27865_ (.A(_02697_),
    .B(_02699_),
    .C1(_02690_),
    .C2(_02700_),
    .ZN(_02701_));
 CLKBUF_X2 _27866_ (.A(_02629_),
    .Z(_02702_));
 AND2_X1 _27867_ (.A1(_02695_),
    .A2(_02702_),
    .ZN(_02703_));
 AND2_X2 _27868_ (.A1(_02674_),
    .A2(_02652_),
    .ZN(_02704_));
 NAND2_X1 _27869_ (.A1(_02695_),
    .A2(_02704_),
    .ZN(_02705_));
 NAND3_X1 _27870_ (.A1(_02675_),
    .A2(_02694_),
    .A3(_02678_),
    .ZN(_02706_));
 NAND2_X1 _27871_ (.A1(_02705_),
    .A2(_02706_),
    .ZN(_02707_));
 NOR4_X1 _27872_ (.A1(_02692_),
    .A2(_02701_),
    .A3(_02703_),
    .A4(_02707_),
    .ZN(_02708_));
 AND2_X1 _27873_ (.A1(_02622_),
    .A2(_02694_),
    .ZN(_02709_));
 AND2_X1 _27874_ (.A1(_02638_),
    .A2(_02656_),
    .ZN(_02710_));
 BUF_X2 _27875_ (.A(_02710_),
    .Z(_02711_));
 NAND2_X1 _27876_ (.A1(_02709_),
    .A2(_02711_),
    .ZN(_02712_));
 INV_X1 _27877_ (.A(_02709_),
    .ZN(_02713_));
 AND2_X1 _27878_ (.A1(_02627_),
    .A2(_02656_),
    .ZN(_02714_));
 INV_X1 _27879_ (.A(_02714_),
    .ZN(_02715_));
 OAI21_X1 _27880_ (.A(_02712_),
    .B1(_02713_),
    .B2(_02715_),
    .ZN(_02716_));
 BUF_X2 _27881_ (.A(_02709_),
    .Z(_02717_));
 AOI21_X1 _27882_ (.A(_02716_),
    .B1(_02647_),
    .B2(_02717_),
    .ZN(_02718_));
 NOR2_X1 _27883_ (.A1(_02630_),
    .A2(_02669_),
    .ZN(_02719_));
 INV_X1 _27884_ (.A(_02719_),
    .ZN(_02720_));
 OAI21_X1 _27885_ (.A(_02717_),
    .B1(_02720_),
    .B2(_02704_),
    .ZN(_02721_));
 AND2_X1 _27886_ (.A1(_02622_),
    .A2(_02676_),
    .ZN(_02722_));
 BUF_X2 _27887_ (.A(_02722_),
    .Z(_02723_));
 AND2_X2 _27888_ (.A1(_02638_),
    .A2(_02666_),
    .ZN(_02724_));
 OAI21_X1 _27889_ (.A(_02723_),
    .B1(_02654_),
    .B2(_02724_),
    .ZN(_02725_));
 AND2_X1 _27890_ (.A1(_02629_),
    .A2(_16776_),
    .ZN(_02726_));
 CLKBUF_X2 _27891_ (.A(_02726_),
    .Z(_02727_));
 AND2_X2 _27892_ (.A1(_02674_),
    .A2(_02626_),
    .ZN(_02728_));
 OAI21_X1 _27893_ (.A(_02723_),
    .B1(_02727_),
    .B2(_02728_),
    .ZN(_02729_));
 AND4_X1 _27894_ (.A1(_02718_),
    .A2(_02721_),
    .A3(_02725_),
    .A4(_02729_),
    .ZN(_02730_));
 AND2_X1 _27895_ (.A1(_02623_),
    .A2(_02677_),
    .ZN(_02731_));
 BUF_X2 _27896_ (.A(_02731_),
    .Z(_02732_));
 BUF_X2 _27897_ (.A(_02732_),
    .Z(_02733_));
 AND2_X1 _27898_ (.A1(_02674_),
    .A2(_02636_),
    .ZN(_02734_));
 OAI21_X1 _27899_ (.A(_02733_),
    .B1(_02727_),
    .B2(_02734_),
    .ZN(_02735_));
 AND2_X1 _27900_ (.A1(_02662_),
    .A2(_02678_),
    .ZN(_02736_));
 AND2_X1 _27901_ (.A1(_02656_),
    .A2(_02642_),
    .ZN(_02737_));
 NAND2_X1 _27902_ (.A1(_02736_),
    .A2(_02737_),
    .ZN(_02738_));
 NAND2_X1 _27903_ (.A1(_02698_),
    .A2(_02736_),
    .ZN(_02739_));
 NAND3_X1 _27904_ (.A1(_02696_),
    .A2(_02662_),
    .A3(_02678_),
    .ZN(_02740_));
 AND3_X1 _27905_ (.A1(_02738_),
    .A2(_02739_),
    .A3(_02740_),
    .ZN(_02741_));
 BUF_X2 _27906_ (.A(_02736_),
    .Z(_02742_));
 INV_X1 _27907_ (.A(_02684_),
    .ZN(_02743_));
 NAND2_X1 _27908_ (.A1(_02743_),
    .A2(_02702_),
    .ZN(_02744_));
 INV_X1 _27909_ (.A(_02744_),
    .ZN(_02745_));
 OAI21_X1 _27910_ (.A(_02742_),
    .B1(_02745_),
    .B2(_02641_),
    .ZN(_02746_));
 BUF_X2 _27911_ (.A(_02626_),
    .Z(_02747_));
 BUF_X2 _27912_ (.A(_02656_),
    .Z(_02748_));
 OAI211_X1 _27913_ (.A(_02732_),
    .B(_02747_),
    .C1(_02667_),
    .C2(_02748_),
    .ZN(_02749_));
 AND4_X1 _27914_ (.A1(_02735_),
    .A2(_02741_),
    .A3(_02746_),
    .A4(_02749_),
    .ZN(_02750_));
 AND4_X1 _27915_ (.A1(_02673_),
    .A2(_02708_),
    .A3(_02730_),
    .A4(_02750_),
    .ZN(_02751_));
 AND2_X1 _27916_ (.A1(_16782_),
    .A2(_16781_),
    .ZN(_02752_));
 AND2_X1 _27917_ (.A1(_02752_),
    .A2(_02623_),
    .ZN(_02753_));
 CLKBUF_X2 _27918_ (.A(_02753_),
    .Z(_02754_));
 AND2_X1 _27919_ (.A1(_02670_),
    .A2(_02754_),
    .ZN(_02755_));
 INV_X1 _27920_ (.A(_02755_),
    .ZN(_02756_));
 AND2_X1 _27921_ (.A1(_02658_),
    .A2(_02754_),
    .ZN(_02757_));
 INV_X1 _27922_ (.A(_02757_),
    .ZN(_02758_));
 BUF_X2 _27923_ (.A(_02754_),
    .Z(_02759_));
 NAND2_X1 _27924_ (.A1(_02759_),
    .A2(_02734_),
    .ZN(_02760_));
 INV_X1 _27925_ (.A(_02652_),
    .ZN(_02761_));
 NAND3_X1 _27926_ (.A1(_02759_),
    .A2(_02761_),
    .A3(_02667_),
    .ZN(_02762_));
 NAND4_X1 _27927_ (.A1(_02756_),
    .A2(_02758_),
    .A3(_02760_),
    .A4(_02762_),
    .ZN(_02763_));
 AND2_X1 _27928_ (.A1(_02662_),
    .A2(_02752_),
    .ZN(_02764_));
 AND2_X2 _27929_ (.A1(_02639_),
    .A2(_02684_),
    .ZN(_02765_));
 AND2_X1 _27930_ (.A1(_02764_),
    .A2(_02765_),
    .ZN(_02766_));
 AND3_X1 _27931_ (.A1(_02704_),
    .A2(_02662_),
    .A3(_02752_),
    .ZN(_02767_));
 OR2_X1 _27932_ (.A1(_02766_),
    .A2(_02767_),
    .ZN(_02768_));
 CLKBUF_X2 _27933_ (.A(_02764_),
    .Z(_02769_));
 OAI211_X1 _27934_ (.A(_02769_),
    .B(_02748_),
    .C1(_02747_),
    .C2(_02642_),
    .ZN(_02770_));
 NAND2_X1 _27935_ (.A1(_02769_),
    .A2(_02696_),
    .ZN(_02771_));
 INV_X1 _27936_ (.A(_02769_),
    .ZN(_02772_));
 INV_X1 _27937_ (.A(_02698_),
    .ZN(_02773_));
 OAI211_X1 _27938_ (.A(_02770_),
    .B(_02771_),
    .C1(_02772_),
    .C2(_02773_),
    .ZN(_02774_));
 INV_X1 _27939_ (.A(_02638_),
    .ZN(_02775_));
 NAND2_X1 _27940_ (.A1(_02775_),
    .A2(_02702_),
    .ZN(_02776_));
 NOR2_X1 _27941_ (.A1(_02772_),
    .A2(_02776_),
    .ZN(_02777_));
 NOR4_X1 _27942_ (.A1(_02763_),
    .A2(_02768_),
    .A3(_02774_),
    .A4(_02777_),
    .ZN(_02778_));
 AND2_X1 _27943_ (.A1(_02694_),
    .A2(_02752_),
    .ZN(_02779_));
 CLKBUF_X2 _27944_ (.A(_02779_),
    .Z(_02780_));
 NAND2_X1 _27945_ (.A1(_02698_),
    .A2(_02780_),
    .ZN(_02781_));
 BUF_X2 _27946_ (.A(_02714_),
    .Z(_02782_));
 NAND2_X1 _27947_ (.A1(_02782_),
    .A2(_02780_),
    .ZN(_02783_));
 AND2_X1 _27948_ (.A1(_02781_),
    .A2(_02783_),
    .ZN(_02784_));
 AND2_X1 _27949_ (.A1(_02752_),
    .A2(_02676_),
    .ZN(_02785_));
 AND2_X1 _27950_ (.A1(_02632_),
    .A2(_02785_),
    .ZN(_02786_));
 INV_X1 _27951_ (.A(_02786_),
    .ZN(_02787_));
 AND2_X1 _27952_ (.A1(_02640_),
    .A2(_02785_),
    .ZN(_02788_));
 INV_X1 _27953_ (.A(_02788_),
    .ZN(_02789_));
 AND2_X1 _27954_ (.A1(_02643_),
    .A2(_02785_),
    .ZN(_02790_));
 INV_X1 _27955_ (.A(_02790_),
    .ZN(_02791_));
 AND3_X1 _27956_ (.A1(_02656_),
    .A2(_02752_),
    .A3(_02676_),
    .ZN(_02792_));
 AND2_X1 _27957_ (.A1(_02684_),
    .A2(_02666_),
    .ZN(_02793_));
 AOI22_X1 _27958_ (.A1(_02792_),
    .A2(_02743_),
    .B1(_02793_),
    .B2(_02785_),
    .ZN(_02794_));
 AND4_X1 _27959_ (.A1(_02787_),
    .A2(_02789_),
    .A3(_02791_),
    .A4(_02794_),
    .ZN(_02795_));
 AND2_X2 _27960_ (.A1(_02629_),
    .A2(_02652_),
    .ZN(_02796_));
 AND2_X1 _27961_ (.A1(_02780_),
    .A2(_02796_),
    .ZN(_02797_));
 INV_X1 _27962_ (.A(_02797_),
    .ZN(_02798_));
 BUF_X2 _27963_ (.A(_02780_),
    .Z(_02799_));
 CLKBUF_X2 _27964_ (.A(_02674_),
    .Z(_02800_));
 OAI211_X1 _27965_ (.A(_02799_),
    .B(_02800_),
    .C1(_02747_),
    .C2(_02657_),
    .ZN(_02801_));
 AND4_X1 _27966_ (.A1(_02784_),
    .A2(_02795_),
    .A3(_02798_),
    .A4(_02801_),
    .ZN(_02802_));
 NOR2_X1 _27967_ (.A1(_02620_),
    .A2(_16781_),
    .ZN(_02803_));
 AND2_X1 _27968_ (.A1(_02803_),
    .A2(_02694_),
    .ZN(_02804_));
 CLKBUF_X2 _27969_ (.A(_02804_),
    .Z(_02805_));
 OAI21_X1 _27970_ (.A(_02805_),
    .B1(_02737_),
    .B2(_02647_),
    .ZN(_02806_));
 INV_X1 _27971_ (.A(_02704_),
    .ZN(_02807_));
 INV_X1 _27972_ (.A(_02765_),
    .ZN(_02808_));
 NAND2_X1 _27973_ (.A1(_02807_),
    .A2(_02808_),
    .ZN(_02809_));
 OAI21_X1 _27974_ (.A(_02805_),
    .B1(_02720_),
    .B2(_02809_),
    .ZN(_02810_));
 AND2_X1 _27975_ (.A1(_02803_),
    .A2(_02676_),
    .ZN(_02811_));
 BUF_X2 _27976_ (.A(_02811_),
    .Z(_02812_));
 CLKBUF_X2 _27977_ (.A(_02632_),
    .Z(_02813_));
 NAND2_X1 _27978_ (.A1(_02812_),
    .A2(_02813_),
    .ZN(_02814_));
 AND2_X1 _27979_ (.A1(_02652_),
    .A2(_02646_),
    .ZN(_02815_));
 INV_X1 _27980_ (.A(_02815_),
    .ZN(_02816_));
 INV_X1 _27981_ (.A(_02793_),
    .ZN(_02817_));
 NAND2_X1 _27982_ (.A1(_02816_),
    .A2(_02817_),
    .ZN(_02818_));
 OAI21_X1 _27983_ (.A(_02811_),
    .B1(_02818_),
    .B2(_02711_),
    .ZN(_02819_));
 AND4_X1 _27984_ (.A1(_02806_),
    .A2(_02810_),
    .A3(_02814_),
    .A4(_02819_),
    .ZN(_02820_));
 AND2_X1 _27985_ (.A1(_02662_),
    .A2(_02803_),
    .ZN(_02821_));
 NAND2_X1 _27986_ (.A1(_02821_),
    .A2(_02793_),
    .ZN(_02822_));
 AND2_X1 _27987_ (.A1(_02803_),
    .A2(_02623_),
    .ZN(_02823_));
 AND2_X1 _27988_ (.A1(_02823_),
    .A2(_02682_),
    .ZN(_02824_));
 INV_X1 _27989_ (.A(_02824_),
    .ZN(_02825_));
 NAND2_X1 _27990_ (.A1(_02726_),
    .A2(_02823_),
    .ZN(_02826_));
 AND2_X1 _27991_ (.A1(_02825_),
    .A2(_02826_),
    .ZN(_02827_));
 BUF_X2 _27992_ (.A(_02821_),
    .Z(_02828_));
 CLKBUF_X2 _27993_ (.A(_02636_),
    .Z(_02829_));
 OAI221_X1 _27994_ (.A(_02828_),
    .B1(_02829_),
    .B2(_02657_),
    .C1(_02800_),
    .C2(_02702_),
    .ZN(_02830_));
 BUF_X2 _27995_ (.A(_02823_),
    .Z(_02831_));
 INV_X1 _27996_ (.A(_02627_),
    .ZN(_02832_));
 AND2_X1 _27997_ (.A1(_02832_),
    .A2(_02656_),
    .ZN(_02833_));
 OAI21_X1 _27998_ (.A(_02831_),
    .B1(_02833_),
    .B2(_02696_),
    .ZN(_02834_));
 AND4_X1 _27999_ (.A1(_02822_),
    .A2(_02827_),
    .A3(_02830_),
    .A4(_02834_),
    .ZN(_02835_));
 AND4_X1 _28000_ (.A1(_02778_),
    .A2(_02802_),
    .A3(_02820_),
    .A4(_02835_),
    .ZN(_02836_));
 NAND2_X4 _28001_ (.A1(_02751_),
    .A2(_02836_),
    .ZN(_02837_));
 XNOR2_X1 _28002_ (.A(_02619_),
    .B(_02837_),
    .ZN(_02838_));
 INV_X1 _28003_ (.A(_17131_),
    .ZN(_02839_));
 XNOR2_X1 _28004_ (.A(_02838_),
    .B(_02839_),
    .ZN(_02840_));
 MUX2_X1 _28005_ (.A(_01836_),
    .B(_02840_),
    .S(_01825_),
    .Z(_00708_));
 XOR2_X1 _28006_ (.A(_17089_),
    .B(_17185_),
    .Z(_02841_));
 XOR2_X1 _28007_ (.A(_01600_),
    .B(_02841_),
    .Z(_02842_));
 XNOR2_X1 _28008_ (.A(_14368_),
    .B(_02842_),
    .ZN(_02843_));
 MUX2_X1 _28009_ (.A(_01252_),
    .B(_02843_),
    .S(_01780_),
    .Z(_01176_));
 XNOR2_X1 _28010_ (.A(_17092_),
    .B(_17188_),
    .ZN(_02844_));
 XNOR2_X1 _28011_ (.A(_01603_),
    .B(_02844_),
    .ZN(_02845_));
 BUF_X2 _28012_ (.A(_03933_),
    .Z(_02846_));
 MUX2_X1 _28013_ (.A(_01263_),
    .B(_02845_),
    .S(_02846_),
    .Z(_01179_));
 XNOR2_X1 _28014_ (.A(_17093_),
    .B(_17189_),
    .ZN(_02847_));
 XNOR2_X1 _28015_ (.A(_01606_),
    .B(_02847_),
    .ZN(_02848_));
 MUX2_X1 _28016_ (.A(_01274_),
    .B(_02848_),
    .S(_02846_),
    .Z(_01180_));
 XOR2_X1 _28017_ (.A(_17094_),
    .B(_17190_),
    .Z(_02849_));
 XOR2_X1 _28018_ (.A(_01607_),
    .B(_02849_),
    .Z(_02850_));
 XNOR2_X1 _28019_ (.A(_14554_),
    .B(_02850_),
    .ZN(_02851_));
 MUX2_X1 _28020_ (.A(_01285_),
    .B(_02851_),
    .S(_02846_),
    .Z(_01181_));
 XNOR2_X1 _28021_ (.A(_17095_),
    .B(_17191_),
    .ZN(_02852_));
 NOR2_X1 _28022_ (.A1(_03933_),
    .A2(_01296_),
    .ZN(_02853_));
 AOI21_X1 _28023_ (.A(_02853_),
    .B1(_02852_),
    .B2(_01736_),
    .ZN(_02854_));
 NAND2_X1 _28024_ (.A1(_01610_),
    .A2(_03738_),
    .ZN(_02855_));
 MUX2_X1 _28025_ (.A(_02852_),
    .B(_02854_),
    .S(_02855_),
    .Z(_01182_));
 XNOR2_X1 _28026_ (.A(_17096_),
    .B(_17192_),
    .ZN(_02856_));
 XNOR2_X1 _28027_ (.A(_01612_),
    .B(_02856_),
    .ZN(_02857_));
 MUX2_X1 _28028_ (.A(_01307_),
    .B(_02857_),
    .S(_02846_),
    .Z(_01183_));
 XNOR2_X1 _28029_ (.A(_10932_),
    .B(_17193_),
    .ZN(_02858_));
 XNOR2_X1 _28030_ (.A(_01614_),
    .B(_02858_),
    .ZN(_02859_));
 MUX2_X1 _28031_ (.A(_01318_),
    .B(_02859_),
    .S(_02846_),
    .Z(_01184_));
 XOR2_X1 _28032_ (.A(_10938_),
    .B(_17194_),
    .Z(_02860_));
 XNOR2_X1 _28033_ (.A(_01617_),
    .B(_02860_),
    .ZN(_02861_));
 MUX2_X1 _28034_ (.A(_01329_),
    .B(_02861_),
    .S(_02846_),
    .Z(_01185_));
 XOR2_X1 _28035_ (.A(_17068_),
    .B(_17164_),
    .Z(_02862_));
 XOR2_X1 _28036_ (.A(_01618_),
    .B(_02862_),
    .Z(_02863_));
 XNOR2_X1 _28037_ (.A(_15064_),
    .B(_02863_),
    .ZN(_02864_));
 MUX2_X1 _28038_ (.A(_01213_),
    .B(_02864_),
    .S(_02846_),
    .Z(_01155_));
 XOR2_X1 _28039_ (.A(_17069_),
    .B(_17165_),
    .Z(_02865_));
 XOR2_X1 _28040_ (.A(_01621_),
    .B(_02865_),
    .Z(_02866_));
 XNOR2_X1 _28041_ (.A(_15145_),
    .B(_02866_),
    .ZN(_02867_));
 MUX2_X1 _28042_ (.A(_01224_),
    .B(_02867_),
    .S(_02846_),
    .Z(_01156_));
 XOR2_X1 _28043_ (.A(_17142_),
    .B(_17024_),
    .Z(_02868_));
 AND3_X1 _28044_ (.A1(_02499_),
    .A2(_02586_),
    .A3(_02389_),
    .ZN(_02869_));
 AND3_X1 _28045_ (.A1(_02398_),
    .A2(_02586_),
    .A3(_02389_),
    .ZN(_02870_));
 AND2_X1 _28046_ (.A1(_02403_),
    .A2(_16727_),
    .ZN(_02871_));
 AOI211_X1 _28047_ (.A(_02869_),
    .B(_02870_),
    .C1(_02391_),
    .C2(_02871_),
    .ZN(_02872_));
 AND2_X1 _28048_ (.A1(_02465_),
    .A2(_02441_),
    .ZN(_02873_));
 INV_X1 _28049_ (.A(_02873_),
    .ZN(_02874_));
 NAND3_X1 _28050_ (.A1(_02526_),
    .A2(_02389_),
    .A3(_02436_),
    .ZN(_02875_));
 NAND3_X1 _28051_ (.A1(_02476_),
    .A2(_02389_),
    .A3(_02436_),
    .ZN(_02876_));
 NAND4_X1 _28052_ (.A1(_02401_),
    .A2(_02413_),
    .A3(_02436_),
    .A4(_02389_),
    .ZN(_02877_));
 AND4_X1 _28053_ (.A1(_02874_),
    .A2(_02875_),
    .A3(_02876_),
    .A4(_02877_),
    .ZN(_02878_));
 NAND2_X1 _28054_ (.A1(_02489_),
    .A2(_02441_),
    .ZN(_02879_));
 BUF_X2 _28055_ (.A(_02399_),
    .Z(_02880_));
 OAI211_X1 _28056_ (.A(_02461_),
    .B(_02394_),
    .C1(_02880_),
    .C2(_02557_),
    .ZN(_02881_));
 OAI21_X1 _28057_ (.A(_02461_),
    .B1(_02595_),
    .B2(_02522_),
    .ZN(_02882_));
 AND4_X1 _28058_ (.A1(_02878_),
    .A2(_02879_),
    .A3(_02881_),
    .A4(_02882_),
    .ZN(_02883_));
 NAND3_X1 _28059_ (.A1(_02527_),
    .A2(_02586_),
    .A3(_02389_),
    .ZN(_02884_));
 INV_X1 _28060_ (.A(_02390_),
    .ZN(_02885_));
 OAI21_X1 _28061_ (.A(_02884_),
    .B1(_02885_),
    .B2(_02589_),
    .ZN(_02886_));
 AND2_X2 _28062_ (.A1(_02401_),
    .A2(_02413_),
    .ZN(_02887_));
 AOI21_X1 _28063_ (.A(_02886_),
    .B1(_02391_),
    .B2(_02887_),
    .ZN(_02888_));
 NAND2_X1 _28064_ (.A1(_02527_),
    .A2(_02432_),
    .ZN(_02889_));
 NAND2_X1 _28065_ (.A1(_02432_),
    .A2(_02522_),
    .ZN(_02890_));
 OAI211_X1 _28066_ (.A(_02889_),
    .B(_02890_),
    .C1(_02425_),
    .C2(_02419_),
    .ZN(_02891_));
 AOI21_X1 _28067_ (.A(_02419_),
    .B1(_02447_),
    .B2(_02444_),
    .ZN(_02892_));
 AND4_X1 _28068_ (.A1(_02429_),
    .A2(_02394_),
    .A3(_02389_),
    .A4(_02558_),
    .ZN(_02893_));
 NOR3_X1 _28069_ (.A1(_02891_),
    .A2(_02892_),
    .A3(_02893_),
    .ZN(_02894_));
 AND4_X1 _28070_ (.A1(_02872_),
    .A2(_02883_),
    .A3(_02888_),
    .A4(_02894_),
    .ZN(_02895_));
 OAI21_X1 _28071_ (.A(_02503_),
    .B1(_02410_),
    .B2(_02467_),
    .ZN(_02896_));
 AND2_X1 _28072_ (.A1(_02394_),
    .A2(_02557_),
    .ZN(_02897_));
 OAI21_X1 _28073_ (.A(_02503_),
    .B1(_02897_),
    .B2(_02570_),
    .ZN(_02898_));
 AND2_X1 _28074_ (.A1(_02896_),
    .A2(_02898_),
    .ZN(_02899_));
 AND2_X1 _28075_ (.A1(_02610_),
    .A2(_02478_),
    .ZN(_02900_));
 INV_X1 _28076_ (.A(_02900_),
    .ZN(_02901_));
 OAI211_X1 _28077_ (.A(_02478_),
    .B(_02434_),
    .C1(_02880_),
    .C2(_02429_),
    .ZN(_02902_));
 OAI211_X1 _28078_ (.A(_02478_),
    .B(_02454_),
    .C1(_02399_),
    .C2(_02557_),
    .ZN(_02903_));
 AND4_X1 _28079_ (.A1(_02487_),
    .A2(_02901_),
    .A3(_02902_),
    .A4(_02903_),
    .ZN(_02904_));
 AND2_X1 _28080_ (.A1(_02508_),
    .A2(_02394_),
    .ZN(_02905_));
 OAI21_X1 _28081_ (.A(_02515_),
    .B1(_02905_),
    .B2(_02551_),
    .ZN(_02906_));
 AND2_X1 _28082_ (.A1(_02905_),
    .A2(_02493_),
    .ZN(_02907_));
 AND2_X1 _28083_ (.A1(_02481_),
    .A2(_02493_),
    .ZN(_02908_));
 AND2_X1 _28084_ (.A1(_02428_),
    .A2(_16730_),
    .ZN(_02909_));
 AND2_X1 _28085_ (.A1(_02492_),
    .A2(_02909_),
    .ZN(_02910_));
 NOR4_X1 _28086_ (.A1(_02907_),
    .A2(_02496_),
    .A3(_02908_),
    .A4(_02910_),
    .ZN(_02911_));
 AND4_X1 _28087_ (.A1(_02899_),
    .A2(_02904_),
    .A3(_02906_),
    .A4(_02911_),
    .ZN(_02912_));
 AND2_X1 _28088_ (.A1(_02905_),
    .A2(_02581_),
    .ZN(_02913_));
 OAI21_X1 _28089_ (.A(_02581_),
    .B1(_02465_),
    .B2(_02467_),
    .ZN(_02914_));
 NAND3_X1 _28090_ (.A1(_02410_),
    .A2(_02417_),
    .A3(_02567_),
    .ZN(_02915_));
 OAI211_X1 _28091_ (.A(_02914_),
    .B(_02915_),
    .C1(_02409_),
    .C2(_02569_),
    .ZN(_02916_));
 AOI211_X1 _28092_ (.A(_02913_),
    .B(_02916_),
    .C1(_02581_),
    .C2(_02871_),
    .ZN(_02917_));
 AND2_X1 _28093_ (.A1(_02593_),
    .A2(_02563_),
    .ZN(_02918_));
 NAND3_X1 _28094_ (.A1(_02602_),
    .A2(_02567_),
    .A3(_02459_),
    .ZN(_02919_));
 OAI211_X1 _28095_ (.A(_02608_),
    .B(_02919_),
    .C1(_02612_),
    .C2(_02544_),
    .ZN(_02920_));
 AND2_X1 _28096_ (.A1(_02519_),
    .A2(_02508_),
    .ZN(_02921_));
 AOI211_X1 _28097_ (.A(_02918_),
    .B(_02920_),
    .C1(_02593_),
    .C2(_02921_),
    .ZN(_02922_));
 NAND2_X1 _28098_ (.A1(_02575_),
    .A2(_02887_),
    .ZN(_02923_));
 AND2_X1 _28099_ (.A1(_02393_),
    .A2(_02423_),
    .ZN(_02924_));
 OAI211_X1 _28100_ (.A(_02586_),
    .B(_02583_),
    .C1(_02924_),
    .C2(_02446_),
    .ZN(_02925_));
 NOR2_X2 _28101_ (.A1(_02427_),
    .A2(_02400_),
    .ZN(_02926_));
 INV_X1 _28102_ (.A(_02397_),
    .ZN(_02927_));
 NAND4_X1 _28103_ (.A1(_02926_),
    .A2(_02586_),
    .A3(_02927_),
    .A4(_02567_),
    .ZN(_02928_));
 NAND2_X1 _28104_ (.A1(_02574_),
    .A2(_02466_),
    .ZN(_02929_));
 AND4_X1 _28105_ (.A1(_02923_),
    .A2(_02925_),
    .A3(_02928_),
    .A4(_02929_),
    .ZN(_02930_));
 AND2_X1 _28106_ (.A1(_02599_),
    .A2(_02486_),
    .ZN(_02931_));
 INV_X1 _28107_ (.A(_02599_),
    .ZN(_02932_));
 INV_X1 _28108_ (.A(_02467_),
    .ZN(_02933_));
 OAI21_X1 _28109_ (.A(_02604_),
    .B1(_02932_),
    .B2(_02933_),
    .ZN(_02934_));
 AOI211_X1 _28110_ (.A(_02931_),
    .B(_02934_),
    .C1(_02599_),
    .C2(_02897_),
    .ZN(_02935_));
 AND4_X1 _28111_ (.A1(_02917_),
    .A2(_02922_),
    .A3(_02930_),
    .A4(_02935_),
    .ZN(_02936_));
 NAND4_X1 _28112_ (.A1(_02532_),
    .A2(_02557_),
    .A3(_02459_),
    .A4(_02403_),
    .ZN(_02937_));
 INV_X2 _28113_ (.A(_02548_),
    .ZN(_02938_));
 OAI21_X1 _28114_ (.A(_02937_),
    .B1(_02490_),
    .B2(_02938_),
    .ZN(_02939_));
 NAND2_X1 _28115_ (.A1(_02408_),
    .A2(_02548_),
    .ZN(_02940_));
 OAI21_X1 _28116_ (.A(_02940_),
    .B1(_02411_),
    .B2(_02938_),
    .ZN(_02941_));
 AND4_X1 _28117_ (.A1(_02429_),
    .A2(_02434_),
    .A3(_02532_),
    .A4(_02459_),
    .ZN(_02942_));
 NOR3_X1 _28118_ (.A1(_02939_),
    .A2(_02941_),
    .A3(_02942_),
    .ZN(_02943_));
 AND2_X1 _28119_ (.A1(_02533_),
    .A2(_02465_),
    .ZN(_02944_));
 NAND2_X1 _28120_ (.A1(_02533_),
    .A2(_02450_),
    .ZN(_02945_));
 NAND3_X1 _28121_ (.A1(_02404_),
    .A2(_02387_),
    .A3(_02532_),
    .ZN(_02946_));
 NAND2_X1 _28122_ (.A1(_02945_),
    .A2(_02946_),
    .ZN(_02947_));
 AOI211_X1 _28123_ (.A(_02944_),
    .B(_02947_),
    .C1(_02454_),
    .C2(_02534_),
    .ZN(_02948_));
 NAND2_X1 _28124_ (.A1(_02547_),
    .A2(_02560_),
    .ZN(_02949_));
 NAND3_X1 _28125_ (.A1(_02519_),
    .A2(_02560_),
    .A3(_02508_),
    .ZN(_02950_));
 NAND4_X1 _28126_ (.A1(_02472_),
    .A2(_02532_),
    .A3(_02403_),
    .A4(_02417_),
    .ZN(_02951_));
 NAND2_X1 _28127_ (.A1(_02560_),
    .A2(_02476_),
    .ZN(_02952_));
 AND4_X1 _28128_ (.A1(_02949_),
    .A2(_02950_),
    .A3(_02951_),
    .A4(_02952_),
    .ZN(_02953_));
 AND2_X1 _28129_ (.A1(_02537_),
    .A2(_02494_),
    .ZN(_02954_));
 INV_X1 _28130_ (.A(_02954_),
    .ZN(_02955_));
 AND2_X1 _28131_ (.A1(_02537_),
    .A2(_02602_),
    .ZN(_02956_));
 INV_X1 _28132_ (.A(_02956_),
    .ZN(_02957_));
 NAND2_X1 _28133_ (.A1(_02398_),
    .A2(_02537_),
    .ZN(_02958_));
 NAND2_X1 _28134_ (.A1(_02605_),
    .A2(_02537_),
    .ZN(_02959_));
 AND4_X1 _28135_ (.A1(_02955_),
    .A2(_02957_),
    .A3(_02958_),
    .A4(_02959_),
    .ZN(_02960_));
 AND4_X1 _28136_ (.A1(_02943_),
    .A2(_02948_),
    .A3(_02953_),
    .A4(_02960_),
    .ZN(_02961_));
 NAND4_X1 _28137_ (.A1(_02895_),
    .A2(_02912_),
    .A3(_02936_),
    .A4(_02961_),
    .ZN(_02962_));
 NOR2_X2 _28138_ (.A1(_02962_),
    .A2(_02616_),
    .ZN(_02963_));
 AND2_X1 _28139_ (.A1(_01901_),
    .A2(_01953_),
    .ZN(_02964_));
 INV_X1 _28140_ (.A(_02964_),
    .ZN(_02965_));
 NAND2_X1 _28141_ (.A1(_01901_),
    .A2(_02108_),
    .ZN(_02966_));
 NAND2_X1 _28142_ (.A1(_02032_),
    .A2(_01901_),
    .ZN(_02967_));
 AND3_X1 _28143_ (.A1(_02965_),
    .A2(_02966_),
    .A3(_02967_),
    .ZN(_02968_));
 AND2_X1 _28144_ (.A1(_01882_),
    .A2(_01901_),
    .ZN(_02969_));
 INV_X1 _28145_ (.A(_02969_),
    .ZN(_02970_));
 INV_X1 _28146_ (.A(_01986_),
    .ZN(_02971_));
 OAI21_X1 _28147_ (.A(_01983_),
    .B1(_02971_),
    .B2(_01868_),
    .ZN(_02972_));
 OAI21_X1 _28148_ (.A(_01983_),
    .B1(_02000_),
    .B2(_01924_),
    .ZN(_02973_));
 NAND4_X1 _28149_ (.A1(_02968_),
    .A2(_02970_),
    .A3(_02972_),
    .A4(_02973_),
    .ZN(_02974_));
 NAND4_X1 _28150_ (.A1(_01894_),
    .A2(_01980_),
    .A3(_02103_),
    .A4(_01875_),
    .ZN(_02975_));
 NAND2_X1 _28151_ (.A1(_01899_),
    .A2(_02975_),
    .ZN(_02976_));
 INV_X1 _28152_ (.A(_01897_),
    .ZN(_02977_));
 INV_X1 _28153_ (.A(_02076_),
    .ZN(_02978_));
 AOI21_X1 _28154_ (.A(_02977_),
    .B1(_02978_),
    .B2(_02077_),
    .ZN(_02979_));
 AND2_X1 _28155_ (.A1(_01960_),
    .A2(_01948_),
    .ZN(_02980_));
 AND2_X1 _28156_ (.A1(_01960_),
    .A2(_01938_),
    .ZN(_02981_));
 AND2_X1 _28157_ (.A1(_01960_),
    .A2(_02036_),
    .ZN(_02982_));
 AND4_X1 _28158_ (.A1(_01854_),
    .A2(_01881_),
    .A3(_01896_),
    .A4(_01845_),
    .ZN(_02983_));
 OR4_X1 _28159_ (.A1(_02980_),
    .A2(_02981_),
    .A3(_02982_),
    .A4(_02983_),
    .ZN(_02984_));
 NOR4_X1 _28160_ (.A1(_02974_),
    .A2(_02976_),
    .A3(_02979_),
    .A4(_02984_),
    .ZN(_02985_));
 AND2_X1 _28161_ (.A1(_02009_),
    .A2(_01850_),
    .ZN(_02986_));
 NAND2_X1 _28162_ (.A1(_02986_),
    .A2(_01958_),
    .ZN(_02987_));
 NAND2_X1 _28163_ (.A1(_01989_),
    .A2(_01958_),
    .ZN(_02988_));
 NAND2_X1 _28164_ (.A1(_01958_),
    .A2(_01938_),
    .ZN(_02989_));
 AND4_X1 _28165_ (.A1(_01977_),
    .A2(_02987_),
    .A3(_02988_),
    .A4(_02989_),
    .ZN(_02990_));
 AND3_X1 _28166_ (.A1(_01910_),
    .A2(_01854_),
    .A3(_01932_),
    .ZN(_02991_));
 NAND2_X1 _28167_ (.A1(_01850_),
    .A2(_01906_),
    .ZN(_02992_));
 OAI21_X1 _28168_ (.A(_02124_),
    .B1(_02125_),
    .B2(_02992_),
    .ZN(_02993_));
 AOI211_X1 _28169_ (.A(_02991_),
    .B(_02993_),
    .C1(_02035_),
    .C2(_01952_),
    .ZN(_02994_));
 OAI21_X1 _28170_ (.A(_01934_),
    .B1(_02986_),
    .B2(_01928_),
    .ZN(_02995_));
 NAND2_X1 _28171_ (.A1(_01915_),
    .A2(_01975_),
    .ZN(_02996_));
 OAI21_X1 _28172_ (.A(_01975_),
    .B1(_01884_),
    .B2(_02007_),
    .ZN(_02997_));
 NAND4_X1 _28173_ (.A1(_01867_),
    .A2(_01861_),
    .A3(_01886_),
    .A4(_01932_),
    .ZN(_02998_));
 OAI211_X1 _28174_ (.A(_01975_),
    .B(_01938_),
    .C1(_01861_),
    .C2(_01920_),
    .ZN(_02999_));
 AND4_X1 _28175_ (.A1(_02996_),
    .A2(_02997_),
    .A3(_02998_),
    .A4(_02999_),
    .ZN(_03000_));
 AND4_X1 _28176_ (.A1(_02990_),
    .A2(_02994_),
    .A3(_02995_),
    .A4(_03000_),
    .ZN(_03001_));
 CLKBUF_X2 _28177_ (.A(_01838_),
    .Z(_03002_));
 CLKBUF_X2 _28178_ (.A(_02094_),
    .Z(_03003_));
 OAI211_X1 _28179_ (.A(_03002_),
    .B(_03003_),
    .C1(_02098_),
    .C2(_01945_),
    .ZN(_03004_));
 NAND4_X1 _28180_ (.A1(_02057_),
    .A2(_01885_),
    .A3(_03003_),
    .A4(_02072_),
    .ZN(_03005_));
 NAND2_X1 _28181_ (.A1(_02014_),
    .A2(_02113_),
    .ZN(_03006_));
 NAND2_X1 _28182_ (.A1(_01855_),
    .A2(_02037_),
    .ZN(_03007_));
 NAND4_X1 _28183_ (.A1(_03004_),
    .A2(_03005_),
    .A3(_03006_),
    .A4(_03007_),
    .ZN(_03008_));
 OAI21_X1 _28184_ (.A(_01842_),
    .B1(_01989_),
    .B2(_01911_),
    .ZN(_03009_));
 OAI21_X1 _28185_ (.A(_01842_),
    .B1(_02108_),
    .B2(_01953_),
    .ZN(_03010_));
 OAI211_X1 _28186_ (.A(_03009_),
    .B(_03010_),
    .C1(_02100_),
    .C2(_02992_),
    .ZN(_03011_));
 NAND3_X1 _28187_ (.A1(_01890_),
    .A2(_02006_),
    .A3(_02009_),
    .ZN(_03012_));
 NAND4_X1 _28188_ (.A1(_01885_),
    .A2(_01851_),
    .A3(_01922_),
    .A4(_01887_),
    .ZN(_03013_));
 NAND4_X1 _28189_ (.A1(_02116_),
    .A2(_03012_),
    .A3(_02112_),
    .A4(_03013_),
    .ZN(_03014_));
 OAI21_X1 _28190_ (.A(_02047_),
    .B1(_02986_),
    .B2(_01847_),
    .ZN(_03015_));
 OAI21_X1 _28191_ (.A(_02047_),
    .B1(_01911_),
    .B2(_01912_),
    .ZN(_03016_));
 NAND3_X1 _28192_ (.A1(_01885_),
    .A2(_01905_),
    .A3(_01875_),
    .ZN(_03017_));
 NAND3_X1 _28193_ (.A1(_03015_),
    .A2(_03016_),
    .A3(_03017_),
    .ZN(_03018_));
 NOR4_X1 _28194_ (.A1(_03008_),
    .A2(_03011_),
    .A3(_03014_),
    .A4(_03018_),
    .ZN(_03019_));
 BUF_X2 _28195_ (.A(_01941_),
    .Z(_03020_));
 NAND3_X1 _28196_ (.A1(_01979_),
    .A2(_02094_),
    .A3(_03020_),
    .ZN(_03021_));
 NAND4_X1 _28197_ (.A1(_02094_),
    .A2(_01867_),
    .A3(_01894_),
    .A4(_03020_),
    .ZN(_03022_));
 INV_X1 _28198_ (.A(_02031_),
    .ZN(_03023_));
 OAI211_X1 _28199_ (.A(_03021_),
    .B(_03022_),
    .C1(_03023_),
    .C2(_02077_),
    .ZN(_03024_));
 NAND3_X1 _28200_ (.A1(_01955_),
    .A2(_02094_),
    .A3(_03020_),
    .ZN(_03025_));
 OAI21_X1 _28201_ (.A(_03025_),
    .B1(_03023_),
    .B2(_01988_),
    .ZN(_03026_));
 AND4_X1 _28202_ (.A1(_01846_),
    .A2(_02094_),
    .A3(_01845_),
    .A4(_03020_),
    .ZN(_03027_));
 NOR3_X1 _28203_ (.A1(_03024_),
    .A2(_03026_),
    .A3(_03027_),
    .ZN(_03028_));
 AOI21_X1 _28204_ (.A(_01971_),
    .B1(_02078_),
    .B2(_02101_),
    .ZN(_03029_));
 AND3_X1 _28205_ (.A1(_01928_),
    .A2(_01995_),
    .A3(_02059_),
    .ZN(_03030_));
 AND4_X1 _28206_ (.A1(_01846_),
    .A2(_01850_),
    .A3(_01941_),
    .A4(_01875_),
    .ZN(_03031_));
 NOR4_X1 _28207_ (.A1(_03029_),
    .A2(_03030_),
    .A3(_02023_),
    .A4(_03031_),
    .ZN(_03032_));
 NAND2_X1 _28208_ (.A1(_02079_),
    .A2(_01943_),
    .ZN(_03033_));
 NAND2_X1 _28209_ (.A1(_02000_),
    .A2(_01943_),
    .ZN(_03034_));
 OAI211_X1 _28210_ (.A(_01943_),
    .B(_01905_),
    .C1(_01861_),
    .C2(_01920_),
    .ZN(_03035_));
 AND3_X1 _28211_ (.A1(_03033_),
    .A2(_03034_),
    .A3(_03035_),
    .ZN(_03036_));
 OAI21_X1 _28212_ (.A(_02018_),
    .B1(_01915_),
    .B2(_01963_),
    .ZN(_03037_));
 OAI211_X1 _28213_ (.A(_02018_),
    .B(_01851_),
    .C1(_01861_),
    .C2(_01920_),
    .ZN(_03038_));
 AND2_X1 _28214_ (.A1(_03037_),
    .A2(_03038_),
    .ZN(_03039_));
 AND4_X1 _28215_ (.A1(_03028_),
    .A2(_03032_),
    .A3(_03036_),
    .A4(_03039_),
    .ZN(_03040_));
 NAND4_X1 _28216_ (.A1(_02985_),
    .A2(_03001_),
    .A3(_03019_),
    .A4(_03040_),
    .ZN(_03041_));
 NOR2_X2 _28217_ (.A1(_03041_),
    .A2(_02045_),
    .ZN(_03042_));
 XNOR2_X2 _28218_ (.A(_02963_),
    .B(_03042_),
    .ZN(_03043_));
 XOR2_X1 _28219_ (.A(_02140_),
    .B(_03043_),
    .Z(_03044_));
 MUX2_X1 _28220_ (.A(_02353_),
    .B(_02162_),
    .S(_02188_),
    .Z(_03045_));
 NAND2_X1 _28221_ (.A1(_03045_),
    .A2(_02152_),
    .ZN(_03046_));
 AND2_X1 _28222_ (.A1(_02251_),
    .A2(_02219_),
    .ZN(_03047_));
 AND2_X1 _28223_ (.A1(_02219_),
    .A2(_02194_),
    .ZN(_03048_));
 NOR2_X1 _28224_ (.A1(_03047_),
    .A2(_03048_),
    .ZN(_03049_));
 AND2_X1 _28225_ (.A1(_02195_),
    .A2(_02238_),
    .ZN(_03050_));
 AND2_X1 _28226_ (.A1(_02199_),
    .A2(_02237_),
    .ZN(_03051_));
 BUF_X2 _28227_ (.A(_02238_),
    .Z(_03052_));
 AOI211_X1 _28228_ (.A(_03050_),
    .B(_03051_),
    .C1(_02159_),
    .C2(_03052_),
    .ZN(_03053_));
 OAI21_X1 _28229_ (.A(_03052_),
    .B1(_02363_),
    .B2(_02164_),
    .ZN(_03054_));
 NAND2_X1 _28230_ (.A1(_02246_),
    .A2(_02220_),
    .ZN(_03055_));
 BUF_X2 _28231_ (.A(_02306_),
    .Z(_03056_));
 NAND2_X1 _28232_ (.A1(_02220_),
    .A2(_03056_),
    .ZN(_03057_));
 NAND2_X1 _28233_ (.A1(_02219_),
    .A2(_02361_),
    .ZN(_03058_));
 AND3_X1 _28234_ (.A1(_03055_),
    .A2(_03057_),
    .A3(_03058_),
    .ZN(_03059_));
 AND4_X1 _28235_ (.A1(_03049_),
    .A2(_03053_),
    .A3(_03054_),
    .A4(_03059_),
    .ZN(_03060_));
 NOR3_X2 _28236_ (.A1(_02166_),
    .A2(_16769_),
    .A3(_02155_),
    .ZN(_03061_));
 AND2_X2 _28237_ (.A1(_03061_),
    .A2(_02174_),
    .ZN(_03062_));
 OAI21_X1 _28238_ (.A(_02152_),
    .B1(_03062_),
    .B2(_02221_),
    .ZN(_03063_));
 AND2_X1 _28239_ (.A1(_02330_),
    .A2(_02275_),
    .ZN(_03064_));
 AND2_X1 _28240_ (.A1(_02334_),
    .A2(_02268_),
    .ZN(_03065_));
 AND2_X1 _28241_ (.A1(_02330_),
    .A2(_02252_),
    .ZN(_03066_));
 AND3_X1 _28242_ (.A1(_02248_),
    .A2(_02260_),
    .A3(_02227_),
    .ZN(_03067_));
 NOR4_X1 _28243_ (.A1(_03064_),
    .A2(_03065_),
    .A3(_03066_),
    .A4(_03067_),
    .ZN(_03068_));
 AND4_X1 _28244_ (.A1(_03046_),
    .A2(_03060_),
    .A3(_03063_),
    .A4(_03068_),
    .ZN(_03069_));
 AND3_X1 _28245_ (.A1(_02351_),
    .A2(_02188_),
    .A3(_02240_),
    .ZN(_03070_));
 NAND3_X1 _28246_ (.A1(_02351_),
    .A2(_02145_),
    .A3(_02240_),
    .ZN(_03071_));
 INV_X1 _28247_ (.A(_02246_),
    .ZN(_03072_));
 OAI21_X1 _28248_ (.A(_03071_),
    .B1(_03072_),
    .B2(_02376_),
    .ZN(_03073_));
 AOI211_X1 _28249_ (.A(_03070_),
    .B(_03073_),
    .C1(_02361_),
    .C2(_02380_),
    .ZN(_03074_));
 BUF_X2 _28250_ (.A(_02271_),
    .Z(_03075_));
 OAI211_X1 _28251_ (.A(_02380_),
    .B(_16770_),
    .C1(_03075_),
    .C2(_16769_),
    .ZN(_03076_));
 AND2_X1 _28252_ (.A1(_02324_),
    .A2(_02378_),
    .ZN(_03077_));
 INV_X1 _28253_ (.A(_03077_),
    .ZN(_03078_));
 NAND2_X1 _28254_ (.A1(_02325_),
    .A2(_02288_),
    .ZN(_03079_));
 BUF_X2 _28255_ (.A(_02301_),
    .Z(_03080_));
 AND2_X1 _28256_ (.A1(_02240_),
    .A2(_03080_),
    .ZN(_03081_));
 OAI21_X1 _28257_ (.A(_02326_),
    .B1(_03081_),
    .B2(_02370_),
    .ZN(_03082_));
 AND3_X1 _28258_ (.A1(_03078_),
    .A2(_03079_),
    .A3(_03082_),
    .ZN(_03083_));
 NAND2_X1 _28259_ (.A1(_02259_),
    .A2(_02184_),
    .ZN(_03084_));
 INV_X1 _28260_ (.A(_03084_),
    .ZN(_03085_));
 OAI21_X1 _28261_ (.A(_02339_),
    .B1(_03085_),
    .B2(_02278_),
    .ZN(_03086_));
 OAI21_X1 _28262_ (.A(_02358_),
    .B1(_02176_),
    .B2(_02336_),
    .ZN(_03087_));
 OAI211_X1 _28263_ (.A(_02358_),
    .B(_02352_),
    .C1(_02375_),
    .C2(_02285_),
    .ZN(_03088_));
 OAI211_X1 _28264_ (.A(_02358_),
    .B(_02275_),
    .C1(_02375_),
    .C2(_03080_),
    .ZN(_03089_));
 AND4_X1 _28265_ (.A1(_03086_),
    .A2(_03087_),
    .A3(_03088_),
    .A4(_03089_),
    .ZN(_03090_));
 AND4_X1 _28266_ (.A1(_03074_),
    .A2(_03076_),
    .A3(_03083_),
    .A4(_03090_),
    .ZN(_03091_));
 AND2_X1 _28267_ (.A1(_02173_),
    .A2(_02252_),
    .ZN(_03092_));
 INV_X1 _28268_ (.A(_02173_),
    .ZN(_03093_));
 INV_X1 _28269_ (.A(_02347_),
    .ZN(_03094_));
 INV_X1 _28270_ (.A(_02345_),
    .ZN(_03095_));
 AOI21_X1 _28271_ (.A(_03093_),
    .B1(_03094_),
    .B2(_03095_),
    .ZN(_03096_));
 AOI21_X1 _28272_ (.A(_03093_),
    .B1(_02357_),
    .B2(_02365_),
    .ZN(_03097_));
 AND2_X1 _28273_ (.A1(_02212_),
    .A2(_02254_),
    .ZN(_03098_));
 OR4_X1 _28274_ (.A1(_03092_),
    .A2(_03096_),
    .A3(_03097_),
    .A4(_03098_),
    .ZN(_03099_));
 AND2_X1 _28275_ (.A1(_02328_),
    .A2(_02287_),
    .ZN(_03100_));
 NOR2_X1 _28276_ (.A1(_03100_),
    .A2(_02316_),
    .ZN(_03101_));
 NAND4_X1 _28277_ (.A1(_02284_),
    .A2(_02285_),
    .A3(_02150_),
    .A4(_02162_),
    .ZN(_03102_));
 OAI21_X1 _28278_ (.A(_02369_),
    .B1(_02252_),
    .B2(_02379_),
    .ZN(_03103_));
 OAI21_X1 _28279_ (.A(_02369_),
    .B1(_02200_),
    .B2(_02288_),
    .ZN(_03104_));
 NAND4_X1 _28280_ (.A1(_03101_),
    .A2(_03102_),
    .A3(_03103_),
    .A4(_03104_),
    .ZN(_03105_));
 AND2_X1 _28281_ (.A1(_02209_),
    .A2(_02272_),
    .ZN(_03106_));
 NOR2_X1 _28282_ (.A1(_02322_),
    .A2(_03106_),
    .ZN(_03107_));
 NAND4_X1 _28283_ (.A1(_02284_),
    .A2(_02226_),
    .A3(_02353_),
    .A4(_03080_),
    .ZN(_03108_));
 NAND4_X1 _28284_ (.A1(_02284_),
    .A2(_02352_),
    .A3(_02226_),
    .A4(_03075_),
    .ZN(_03109_));
 NAND4_X1 _28285_ (.A1(_03107_),
    .A2(_02343_),
    .A3(_03108_),
    .A4(_03109_),
    .ZN(_03110_));
 OAI21_X1 _28286_ (.A(_02192_),
    .B1(_02311_),
    .B2(_02337_),
    .ZN(_03111_));
 OAI21_X1 _28287_ (.A(_02191_),
    .B1(_02199_),
    .B2(_02332_),
    .ZN(_03112_));
 INV_X1 _28288_ (.A(_03062_),
    .ZN(_03113_));
 INV_X1 _28289_ (.A(_02191_),
    .ZN(_03114_));
 OAI211_X1 _28290_ (.A(_03111_),
    .B(_03112_),
    .C1(_03113_),
    .C2(_03114_),
    .ZN(_03115_));
 NOR4_X1 _28291_ (.A1(_03099_),
    .A2(_03105_),
    .A3(_03110_),
    .A4(_03115_),
    .ZN(_03116_));
 INV_X1 _28292_ (.A(_02317_),
    .ZN(_03117_));
 NAND2_X1 _28293_ (.A1(_03117_),
    .A2(_03094_),
    .ZN(_03118_));
 OAI21_X1 _28294_ (.A(_02265_),
    .B1(_03118_),
    .B2(_02336_),
    .ZN(_03119_));
 AND2_X1 _28295_ (.A1(_02194_),
    .A2(_02264_),
    .ZN(_03120_));
 INV_X1 _28296_ (.A(_03120_),
    .ZN(_03121_));
 OAI211_X1 _28297_ (.A(_02265_),
    .B(_02275_),
    .C1(_03075_),
    .C2(_03080_),
    .ZN(_03122_));
 AND3_X1 _28298_ (.A1(_03119_),
    .A2(_03121_),
    .A3(_03122_),
    .ZN(_03123_));
 AND2_X1 _28299_ (.A1(_02194_),
    .A2(_02308_),
    .ZN(_03124_));
 AND2_X1 _28300_ (.A1(_02363_),
    .A2(_02274_),
    .ZN(_03125_));
 AND2_X1 _28301_ (.A1(_02268_),
    .A2(_02270_),
    .ZN(_03126_));
 AND2_X1 _28302_ (.A1(_02308_),
    .A2(_02333_),
    .ZN(_03127_));
 NOR4_X1 _28303_ (.A1(_03124_),
    .A2(_03125_),
    .A3(_03126_),
    .A4(_03127_),
    .ZN(_03128_));
 OAI21_X1 _28304_ (.A(_02245_),
    .B1(_02337_),
    .B2(_02327_),
    .ZN(_03129_));
 OAI211_X1 _28305_ (.A(_02260_),
    .B(_02261_),
    .C1(_02221_),
    .C2(_02356_),
    .ZN(_03130_));
 AND3_X1 _28306_ (.A1(_03129_),
    .A2(_03130_),
    .A3(_02255_),
    .ZN(_03131_));
 OAI21_X1 _28307_ (.A(_02235_),
    .B1(_02252_),
    .B2(_02254_),
    .ZN(_03132_));
 NAND2_X1 _28308_ (.A1(_02363_),
    .A2(_02234_),
    .ZN(_03133_));
 NAND3_X1 _28309_ (.A1(_02221_),
    .A2(_02226_),
    .A3(_02261_),
    .ZN(_03134_));
 NAND3_X1 _28310_ (.A1(_02235_),
    .A2(_03080_),
    .A3(_02223_),
    .ZN(_03135_));
 AND4_X1 _28311_ (.A1(_03132_),
    .A2(_03133_),
    .A3(_03134_),
    .A4(_03135_),
    .ZN(_03136_));
 AND4_X1 _28312_ (.A1(_03123_),
    .A2(_03128_),
    .A3(_03131_),
    .A4(_03136_),
    .ZN(_03137_));
 NAND4_X1 _28313_ (.A1(_03069_),
    .A2(_03091_),
    .A3(_03116_),
    .A4(_03137_),
    .ZN(_03138_));
 NOR2_X2 _28314_ (.A1(_03138_),
    .A2(_02282_),
    .ZN(_03139_));
 XNOR2_X1 _28315_ (.A(_03044_),
    .B(_03139_),
    .ZN(_03140_));
 AND2_X1 _28316_ (.A1(_02709_),
    .A2(_02737_),
    .ZN(_03141_));
 INV_X1 _28317_ (.A(_03141_),
    .ZN(_03142_));
 AND2_X1 _28318_ (.A1(_02675_),
    .A2(_02732_),
    .ZN(_03143_));
 INV_X1 _28319_ (.A(_03143_),
    .ZN(_03144_));
 INV_X1 _28320_ (.A(_02696_),
    .ZN(_03145_));
 INV_X1 _28321_ (.A(_02723_),
    .ZN(_03146_));
 OAI211_X1 _28322_ (.A(_03142_),
    .B(_03144_),
    .C1(_03145_),
    .C2(_03146_),
    .ZN(_03147_));
 XNOR2_X2 _28323_ (.A(_02626_),
    .B(_02642_),
    .ZN(_03148_));
 INV_X1 _28324_ (.A(_02674_),
    .ZN(_03149_));
 NOR2_X1 _28325_ (.A1(_03148_),
    .A2(_03149_),
    .ZN(_03150_));
 INV_X1 _28326_ (.A(_03150_),
    .ZN(_03151_));
 INV_X1 _28327_ (.A(_02727_),
    .ZN(_03152_));
 AOI21_X1 _28328_ (.A(_02691_),
    .B1(_03151_),
    .B2(_03152_),
    .ZN(_03153_));
 AND2_X1 _28329_ (.A1(_02703_),
    .A2(_03148_),
    .ZN(_03154_));
 NOR2_X1 _28330_ (.A1(_02782_),
    .A2(_02710_),
    .ZN(_03155_));
 AND2_X1 _28331_ (.A1(_02666_),
    .A2(_02642_),
    .ZN(_03156_));
 INV_X1 _28332_ (.A(_03156_),
    .ZN(_03157_));
 AOI21_X1 _28333_ (.A(_02700_),
    .B1(_03155_),
    .B2(_03157_),
    .ZN(_03158_));
 NOR4_X1 _28334_ (.A1(_03147_),
    .A2(_03153_),
    .A3(_03154_),
    .A4(_03158_),
    .ZN(_03159_));
 INV_X1 _28335_ (.A(_03155_),
    .ZN(_03160_));
 OAI21_X1 _28336_ (.A(_02742_),
    .B1(_03160_),
    .B2(_02671_),
    .ZN(_03161_));
 AND2_X1 _28337_ (.A1(_02739_),
    .A2(_02740_),
    .ZN(_03162_));
 INV_X1 _28338_ (.A(_03162_),
    .ZN(_03163_));
 AND2_X1 _28339_ (.A1(_02724_),
    .A2(_02753_),
    .ZN(_03164_));
 AND3_X1 _28340_ (.A1(_02785_),
    .A2(_02800_),
    .A3(_02627_),
    .ZN(_03165_));
 AND3_X1 _28341_ (.A1(_02753_),
    .A2(_02643_),
    .A3(_02636_),
    .ZN(_03166_));
 NOR4_X1 _28342_ (.A1(_03163_),
    .A2(_03164_),
    .A3(_03165_),
    .A4(_03166_),
    .ZN(_03167_));
 NAND2_X1 _28343_ (.A1(_02743_),
    .A2(_02666_),
    .ZN(_03168_));
 INV_X1 _28344_ (.A(_03168_),
    .ZN(_03169_));
 NAND2_X1 _28345_ (.A1(_03169_),
    .A2(_02733_),
    .ZN(_03170_));
 INV_X1 _28346_ (.A(_02776_),
    .ZN(_03171_));
 BUF_X2 _28347_ (.A(_02764_),
    .Z(_03172_));
 AOI22_X1 _28348_ (.A1(_03171_),
    .A2(_03172_),
    .B1(_02833_),
    .B2(_02831_),
    .ZN(_03173_));
 AND4_X1 _28349_ (.A1(_03161_),
    .A2(_03167_),
    .A3(_03170_),
    .A4(_03173_),
    .ZN(_03174_));
 CLKBUF_X2 _28350_ (.A(_02680_),
    .Z(_03175_));
 OAI21_X1 _28351_ (.A(_03175_),
    .B1(_02670_),
    .B2(_02711_),
    .ZN(_03176_));
 NAND2_X1 _28352_ (.A1(_02686_),
    .A2(_02754_),
    .ZN(_03177_));
 OAI211_X1 _28353_ (.A(_02680_),
    .B(_02642_),
    .C1(_02666_),
    .C2(_02748_),
    .ZN(_03178_));
 AND4_X1 _28354_ (.A1(_02781_),
    .A2(_02649_),
    .A3(_03177_),
    .A4(_03178_),
    .ZN(_03179_));
 AND2_X1 _28355_ (.A1(_02736_),
    .A2(_02765_),
    .ZN(_03180_));
 INV_X1 _28356_ (.A(_03180_),
    .ZN(_03181_));
 AND2_X1 _28357_ (.A1(_02629_),
    .A2(_02684_),
    .ZN(_03182_));
 NAND2_X1 _28358_ (.A1(_03182_),
    .A2(_02732_),
    .ZN(_03183_));
 AOI22_X1 _28359_ (.A1(_02722_),
    .A2(_02686_),
    .B1(_02704_),
    .B2(_02732_),
    .ZN(_03184_));
 NAND3_X1 _28360_ (.A1(_02732_),
    .A2(_02627_),
    .A3(_02748_),
    .ZN(_03185_));
 NAND3_X1 _28361_ (.A1(_02664_),
    .A2(_02829_),
    .A3(_02643_),
    .ZN(_03186_));
 AND4_X1 _28362_ (.A1(_03183_),
    .A2(_03184_),
    .A3(_03185_),
    .A4(_03186_),
    .ZN(_03187_));
 AND4_X1 _28363_ (.A1(_03176_),
    .A2(_03179_),
    .A3(_03181_),
    .A4(_03187_),
    .ZN(_03188_));
 INV_X2 _28364_ (.A(_02823_),
    .ZN(_03189_));
 INV_X1 _28365_ (.A(_02785_),
    .ZN(_03190_));
 OAI22_X1 _28366_ (.A1(_02808_),
    .A2(_03189_),
    .B1(_02773_),
    .B2(_03190_),
    .ZN(_03191_));
 NAND2_X1 _28367_ (.A1(_02635_),
    .A2(_02793_),
    .ZN(_03192_));
 INV_X1 _28368_ (.A(_02821_),
    .ZN(_03193_));
 OAI21_X1 _28369_ (.A(_03192_),
    .B1(_03193_),
    .B2(_02687_),
    .ZN(_03194_));
 AOI211_X1 _28370_ (.A(_03191_),
    .B(_03194_),
    .C1(_02742_),
    .C2(_02745_),
    .ZN(_03195_));
 AND4_X1 _28371_ (.A1(_03159_),
    .A2(_03174_),
    .A3(_03188_),
    .A4(_03195_),
    .ZN(_03196_));
 AOI21_X1 _28372_ (.A(_16778_),
    .B1(_02684_),
    .B2(_02650_),
    .ZN(_03197_));
 NAND3_X1 _28373_ (.A1(_02676_),
    .A2(_02678_),
    .A3(_02628_),
    .ZN(_03198_));
 NOR2_X1 _28374_ (.A1(_03197_),
    .A2(_03198_),
    .ZN(_03199_));
 INV_X1 _28375_ (.A(_02804_),
    .ZN(_03200_));
 NAND3_X1 _28376_ (.A1(_02761_),
    .A2(_02743_),
    .A3(_02666_),
    .ZN(_03201_));
 NOR2_X1 _28377_ (.A1(_03200_),
    .A2(_03201_),
    .ZN(_03202_));
 AND2_X1 _28378_ (.A1(_02629_),
    .A2(_02626_),
    .ZN(_03203_));
 BUF_X2 _28379_ (.A(_02785_),
    .Z(_03204_));
 AOI211_X1 _28380_ (.A(_03199_),
    .B(_03202_),
    .C1(_03203_),
    .C2(_03204_),
    .ZN(_03205_));
 INV_X1 _28381_ (.A(_02780_),
    .ZN(_03206_));
 INV_X1 _28382_ (.A(_02632_),
    .ZN(_03207_));
 AOI21_X1 _28383_ (.A(_03206_),
    .B1(_03152_),
    .B2(_03207_),
    .ZN(_03208_));
 AND2_X2 _28384_ (.A1(_02656_),
    .A2(_02626_),
    .ZN(_03209_));
 NAND2_X1 _28385_ (.A1(_02635_),
    .A2(_03209_),
    .ZN(_03210_));
 CLKBUF_X2 _28386_ (.A(_02803_),
    .Z(_03211_));
 NAND3_X1 _28387_ (.A1(_02671_),
    .A2(_03211_),
    .A3(_02694_),
    .ZN(_03212_));
 NAND2_X1 _28388_ (.A1(_03210_),
    .A2(_03212_),
    .ZN(_03213_));
 AND2_X1 _28389_ (.A1(_02769_),
    .A2(_02658_),
    .ZN(_03214_));
 AND2_X1 _28390_ (.A1(_02675_),
    .A2(_02785_),
    .ZN(_03215_));
 NOR4_X1 _28391_ (.A1(_03208_),
    .A2(_03213_),
    .A3(_03214_),
    .A4(_03215_),
    .ZN(_03216_));
 OAI21_X1 _28392_ (.A(_03172_),
    .B1(_02818_),
    .B2(_02728_),
    .ZN(_03217_));
 OAI21_X1 _28393_ (.A(_02722_),
    .B1(_02682_),
    .B2(_02675_),
    .ZN(_03218_));
 NAND4_X1 _28394_ (.A1(_02622_),
    .A2(_02626_),
    .A3(_02702_),
    .A4(_02676_),
    .ZN(_03219_));
 NAND2_X1 _28395_ (.A1(_03218_),
    .A2(_03219_),
    .ZN(_03220_));
 AND2_X1 _28396_ (.A1(_02727_),
    .A2(_02754_),
    .ZN(_03221_));
 NOR2_X1 _28397_ (.A1(_03220_),
    .A2(_03221_),
    .ZN(_03222_));
 NAND4_X1 _28398_ (.A1(_03205_),
    .A2(_03216_),
    .A3(_03217_),
    .A4(_03222_),
    .ZN(_03223_));
 OAI21_X1 _28399_ (.A(_02828_),
    .B1(_02704_),
    .B2(_02675_),
    .ZN(_03224_));
 NAND2_X1 _28400_ (.A1(_02670_),
    .A2(_02828_),
    .ZN(_03225_));
 AND2_X1 _28401_ (.A1(_03224_),
    .A2(_03225_),
    .ZN(_03226_));
 OAI21_X1 _28402_ (.A(_02799_),
    .B1(_03150_),
    .B2(_02711_),
    .ZN(_03227_));
 OAI21_X1 _28403_ (.A(_02759_),
    .B1(_02813_),
    .B2(_03156_),
    .ZN(_03228_));
 NAND2_X1 _28404_ (.A1(_02775_),
    .A2(_02666_),
    .ZN(_03229_));
 INV_X1 _28405_ (.A(_03229_),
    .ZN(_03230_));
 NAND2_X1 _28406_ (.A1(_03230_),
    .A2(_02831_),
    .ZN(_03231_));
 NAND4_X1 _28407_ (.A1(_03226_),
    .A2(_03227_),
    .A3(_03228_),
    .A4(_03231_),
    .ZN(_03232_));
 NAND2_X1 _28408_ (.A1(_03150_),
    .A2(_02635_),
    .ZN(_03233_));
 BUF_X2 _28409_ (.A(_02623_),
    .Z(_03234_));
 NAND3_X1 _28410_ (.A1(_02796_),
    .A2(_03234_),
    .A3(_02622_),
    .ZN(_03235_));
 AND2_X1 _28411_ (.A1(_03233_),
    .A2(_03235_),
    .ZN(_03236_));
 AND2_X1 _28412_ (.A1(_02666_),
    .A2(_02829_),
    .ZN(_03237_));
 OAI21_X1 _28413_ (.A(_02812_),
    .B1(_03203_),
    .B2(_03237_),
    .ZN(_03238_));
 NAND2_X1 _28414_ (.A1(_02743_),
    .A2(_02800_),
    .ZN(_03239_));
 INV_X1 _28415_ (.A(_03239_),
    .ZN(_03240_));
 AND2_X1 _28416_ (.A1(_03240_),
    .A2(_02811_),
    .ZN(_03241_));
 INV_X1 _28417_ (.A(_03241_),
    .ZN(_03242_));
 NAND2_X1 _28418_ (.A1(_02833_),
    .A2(_02812_),
    .ZN(_03243_));
 NAND4_X1 _28419_ (.A1(_03236_),
    .A2(_03238_),
    .A3(_03242_),
    .A4(_03243_),
    .ZN(_03244_));
 OAI21_X1 _28420_ (.A(_02717_),
    .B1(_03203_),
    .B2(_02704_),
    .ZN(_03245_));
 BUF_X2 _28421_ (.A(_02748_),
    .Z(_03246_));
 OAI21_X1 _28422_ (.A(_02665_),
    .B1(_02647_),
    .B2(_03246_),
    .ZN(_03247_));
 NAND3_X1 _28423_ (.A1(_02709_),
    .A2(_02667_),
    .A3(_02832_),
    .ZN(_03248_));
 NAND3_X1 _28424_ (.A1(_02664_),
    .A2(_02832_),
    .A3(_02702_),
    .ZN(_03249_));
 NAND4_X1 _28425_ (.A1(_03245_),
    .A2(_03247_),
    .A3(_03248_),
    .A4(_03249_),
    .ZN(_03250_));
 NOR4_X1 _28426_ (.A1(_03223_),
    .A2(_03232_),
    .A3(_03244_),
    .A4(_03250_),
    .ZN(_03251_));
 NAND2_X2 _28427_ (.A1(_03196_),
    .A2(_03251_),
    .ZN(_03252_));
 XOR2_X2 _28428_ (.A(_03252_),
    .B(_02837_),
    .Z(_03253_));
 XNOR2_X1 _28429_ (.A(_03140_),
    .B(_03253_),
    .ZN(_03254_));
 XNOR2_X1 _28430_ (.A(_03254_),
    .B(_17142_),
    .ZN(_03255_));
 MUX2_X1 _28431_ (.A(_02868_),
    .B(_03255_),
    .S(_01825_),
    .Z(_00709_));
 XOR2_X1 _28432_ (.A(_17070_),
    .B(_17166_),
    .Z(_03256_));
 XOR2_X1 _28433_ (.A(_01623_),
    .B(_03256_),
    .Z(_03257_));
 XNOR2_X1 _28434_ (.A(_15212_),
    .B(_03257_),
    .ZN(_03258_));
 MUX2_X1 _28435_ (.A(_01233_),
    .B(_03258_),
    .S(_02846_),
    .Z(_01157_));
 XOR2_X1 _28436_ (.A(_17071_),
    .B(_17167_),
    .Z(_03259_));
 XOR2_X1 _28437_ (.A(_01625_),
    .B(_03259_),
    .Z(_03260_));
 XNOR2_X1 _28438_ (.A(_15283_),
    .B(_03260_),
    .ZN(_03261_));
 MUX2_X1 _28439_ (.A(_01234_),
    .B(_03261_),
    .S(_02846_),
    .Z(_01158_));
 XOR2_X1 _28440_ (.A(_17072_),
    .B(_17168_),
    .Z(_03262_));
 XOR2_X1 _28441_ (.A(_01627_),
    .B(_03262_),
    .Z(_03263_));
 XNOR2_X1 _28442_ (.A(_15345_),
    .B(_03263_),
    .ZN(_03264_));
 BUF_X2 _28443_ (.A(_03933_),
    .Z(_03265_));
 MUX2_X1 _28444_ (.A(_01235_),
    .B(_03264_),
    .S(_03265_),
    .Z(_01159_));
 XOR2_X1 _28445_ (.A(_17073_),
    .B(_17169_),
    .Z(_03266_));
 XOR2_X1 _28446_ (.A(_01629_),
    .B(_03266_),
    .Z(_03267_));
 XNOR2_X1 _28447_ (.A(_15405_),
    .B(_03267_),
    .ZN(_03268_));
 MUX2_X1 _28448_ (.A(_01236_),
    .B(_03268_),
    .S(_03265_),
    .Z(_01160_));
 XOR2_X1 _28449_ (.A(_10987_),
    .B(_17138_),
    .Z(_03269_));
 XNOR2_X1 _28450_ (.A(_01761_),
    .B(_03269_),
    .ZN(_03270_));
 XOR2_X1 _28451_ (.A(_15642_),
    .B(_03270_),
    .Z(_03271_));
 MUX2_X1 _28452_ (.A(_01237_),
    .B(_03271_),
    .S(_03265_),
    .Z(_01161_));
 XNOR2_X1 _28453_ (.A(_17107_),
    .B(_17171_),
    .ZN(_03272_));
 XNOR2_X1 _28454_ (.A(_10993_),
    .B(_17139_),
    .ZN(_03273_));
 XOR2_X1 _28455_ (.A(_03272_),
    .B(_03273_),
    .Z(_03274_));
 XNOR2_X1 _28456_ (.A(_15748_),
    .B(_03274_),
    .ZN(_03275_));
 MUX2_X1 _28457_ (.A(_01238_),
    .B(_03275_),
    .S(_03265_),
    .Z(_01162_));
 XOR2_X1 _28458_ (.A(_17076_),
    .B(_17140_),
    .Z(_03276_));
 XNOR2_X1 _28459_ (.A(_01765_),
    .B(_03276_),
    .ZN(_03277_));
 XOR2_X1 _28460_ (.A(_15832_),
    .B(_03277_),
    .Z(_03278_));
 MUX2_X1 _28461_ (.A(_01239_),
    .B(_03278_),
    .S(_03265_),
    .Z(_01163_));
 XOR2_X1 _28462_ (.A(_17077_),
    .B(_17141_),
    .Z(_03279_));
 XOR2_X1 _28463_ (.A(_01768_),
    .B(_03279_),
    .Z(_03280_));
 XNOR2_X1 _28464_ (.A(_15911_),
    .B(_03280_),
    .ZN(_03281_));
 MUX2_X1 _28465_ (.A(_01240_),
    .B(_03281_),
    .S(_03265_),
    .Z(_01164_));
 XOR2_X1 _28466_ (.A(_17111_),
    .B(_17175_),
    .Z(_03282_));
 XOR2_X1 _28467_ (.A(_17079_),
    .B(_17143_),
    .Z(_03283_));
 XNOR2_X1 _28468_ (.A(_03282_),
    .B(_03283_),
    .ZN(_03284_));
 XOR2_X1 _28469_ (.A(_15974_),
    .B(_03284_),
    .Z(_03285_));
 MUX2_X1 _28470_ (.A(_01242_),
    .B(_03285_),
    .S(_03265_),
    .Z(_01166_));
 XOR2_X1 _28471_ (.A(_17112_),
    .B(_17176_),
    .Z(_03286_));
 XOR2_X1 _28472_ (.A(_17080_),
    .B(_17144_),
    .Z(_03287_));
 XNOR2_X1 _28473_ (.A(_03286_),
    .B(_03287_),
    .ZN(_03288_));
 XOR2_X1 _28474_ (.A(_16038_),
    .B(_03288_),
    .Z(_03289_));
 MUX2_X1 _28475_ (.A(_01243_),
    .B(_03289_),
    .S(_03265_),
    .Z(_01167_));
 XOR2_X1 _28476_ (.A(_17153_),
    .B(_17025_),
    .Z(_03290_));
 AND2_X1 _28477_ (.A1(_02391_),
    .A2(_02522_),
    .ZN(_03291_));
 INV_X1 _28478_ (.A(_03291_),
    .ZN(_03292_));
 INV_X1 _28479_ (.A(_02921_),
    .ZN(_03293_));
 OAI211_X1 _28480_ (.A(_03292_),
    .B(_02884_),
    .C1(_03293_),
    .C2(_02885_),
    .ZN(_03294_));
 BUF_X2 _28481_ (.A(_02387_),
    .Z(_03295_));
 NAND3_X1 _28482_ (.A1(_02602_),
    .A2(_03295_),
    .A3(_02438_),
    .ZN(_03296_));
 INV_X1 _28483_ (.A(_02495_),
    .ZN(_03297_));
 OAI21_X1 _28484_ (.A(_03296_),
    .B1(_02885_),
    .B2(_03297_),
    .ZN(_03298_));
 OR3_X1 _28485_ (.A1(_03294_),
    .A2(_02869_),
    .A3(_03298_),
    .ZN(_03299_));
 AOI21_X1 _28486_ (.A(_02419_),
    .B1(_02546_),
    .B2(_03297_),
    .ZN(_03300_));
 OAI211_X1 _28487_ (.A(_02432_),
    .B(_02435_),
    .C1(_02428_),
    .C2(_02430_),
    .ZN(_03301_));
 NAND2_X1 _28488_ (.A1(_02408_),
    .A2(_02418_),
    .ZN(_03302_));
 NAND2_X1 _28489_ (.A1(_03301_),
    .A2(_03302_),
    .ZN(_03303_));
 NOR3_X1 _28490_ (.A1(_03299_),
    .A2(_03300_),
    .A3(_03303_),
    .ZN(_03304_));
 INV_X1 _28491_ (.A(_02450_),
    .ZN(_03305_));
 AOI21_X1 _28492_ (.A(_02938_),
    .B1(_02490_),
    .B2(_03305_),
    .ZN(_03306_));
 INV_X1 _28493_ (.A(_02887_),
    .ZN(_03307_));
 INV_X1 _28494_ (.A(_02466_),
    .ZN(_03308_));
 AOI21_X1 _28495_ (.A(_02938_),
    .B1(_03307_),
    .B2(_03308_),
    .ZN(_03309_));
 AND4_X1 _28496_ (.A1(_02557_),
    .A2(_02553_),
    .A3(_02454_),
    .A4(_02459_),
    .ZN(_03310_));
 OR4_X1 _28497_ (.A1(_02552_),
    .A2(_03306_),
    .A3(_03309_),
    .A4(_03310_),
    .ZN(_03311_));
 OAI21_X1 _28498_ (.A(_02561_),
    .B1(_02500_),
    .B2(_02450_),
    .ZN(_03312_));
 OAI211_X1 _28499_ (.A(_02561_),
    .B(_16730_),
    .C1(_02880_),
    .C2(_02392_),
    .ZN(_03313_));
 OAI21_X1 _28500_ (.A(_02560_),
    .B1(_02578_),
    .B2(_02571_),
    .ZN(_03314_));
 NAND3_X1 _28501_ (.A1(_03312_),
    .A2(_03313_),
    .A3(_03314_),
    .ZN(_03315_));
 OAI21_X1 _28502_ (.A(_02534_),
    .B1(_02466_),
    .B2(_02595_),
    .ZN(_03316_));
 NAND3_X1 _28503_ (.A1(_02541_),
    .A2(_03295_),
    .A3(_02553_),
    .ZN(_03317_));
 NAND2_X1 _28504_ (.A1(_02533_),
    .A2(_02495_),
    .ZN(_03318_));
 NAND3_X1 _28505_ (.A1(_03316_),
    .A2(_03317_),
    .A3(_03318_),
    .ZN(_03319_));
 AND2_X1 _28506_ (.A1(_02887_),
    .A2(_02537_),
    .ZN(_03320_));
 INV_X1 _28507_ (.A(_03320_),
    .ZN(_03321_));
 BUF_X2 _28508_ (.A(_02394_),
    .Z(_03322_));
 OAI211_X1 _28509_ (.A(_02540_),
    .B(_03322_),
    .C1(_02428_),
    .C2(_02430_),
    .ZN(_03323_));
 AND2_X1 _28510_ (.A1(_02511_),
    .A2(_02506_),
    .ZN(_03324_));
 INV_X1 _28511_ (.A(_03324_),
    .ZN(_03325_));
 OAI211_X1 _28512_ (.A(_03321_),
    .B(_03323_),
    .C1(_03325_),
    .C2(_02543_),
    .ZN(_03326_));
 NOR4_X1 _28513_ (.A1(_03311_),
    .A2(_03315_),
    .A3(_03319_),
    .A4(_03326_),
    .ZN(_03327_));
 NAND3_X1 _28514_ (.A1(_02519_),
    .A2(_02442_),
    .A3(_02508_),
    .ZN(_03328_));
 NAND2_X1 _28515_ (.A1(_02926_),
    .A2(_02442_),
    .ZN(_03329_));
 NAND2_X1 _28516_ (.A1(_02500_),
    .A2(_02442_),
    .ZN(_03330_));
 AND3_X1 _28517_ (.A1(_03328_),
    .A2(_03329_),
    .A3(_03330_),
    .ZN(_03331_));
 AND2_X1 _28518_ (.A1(_02450_),
    .A2(_02460_),
    .ZN(_03332_));
 INV_X1 _28519_ (.A(_03332_),
    .ZN(_03333_));
 OAI21_X1 _28520_ (.A(_02462_),
    .B1(_02468_),
    .B2(_02455_),
    .ZN(_03334_));
 NOR2_X1 _28521_ (.A1(_02485_),
    .A2(_02472_),
    .ZN(_03335_));
 NAND3_X1 _28522_ (.A1(_03335_),
    .A2(_02462_),
    .A3(_02927_),
    .ZN(_03336_));
 AND3_X1 _28523_ (.A1(_03333_),
    .A2(_03334_),
    .A3(_03336_),
    .ZN(_03337_));
 NAND4_X1 _28524_ (.A1(_03304_),
    .A2(_03327_),
    .A3(_03331_),
    .A4(_03337_),
    .ZN(_03338_));
 OAI21_X1 _28525_ (.A(_02479_),
    .B1(_02509_),
    .B2(_02571_),
    .ZN(_03339_));
 AOI21_X1 _28526_ (.A(_02516_),
    .B1(_03307_),
    .B2(_03308_),
    .ZN(_03340_));
 AOI21_X1 _28527_ (.A(_03340_),
    .B1(_02476_),
    .B2(_02515_),
    .ZN(_03341_));
 OAI21_X1 _28528_ (.A(_02479_),
    .B1(_02483_),
    .B2(_02455_),
    .ZN(_03342_));
 OAI21_X1 _28529_ (.A(_02515_),
    .B1(_03335_),
    .B2(_03322_),
    .ZN(_03343_));
 AND4_X1 _28530_ (.A1(_03339_),
    .A2(_03341_),
    .A3(_03342_),
    .A4(_03343_),
    .ZN(_03344_));
 NAND2_X1 _28531_ (.A1(_02608_),
    .A2(_02611_),
    .ZN(_03345_));
 INV_X1 _28532_ (.A(_03345_),
    .ZN(_03346_));
 OAI21_X1 _28533_ (.A(_02600_),
    .B1(_02502_),
    .B2(_03324_),
    .ZN(_03347_));
 OAI21_X1 _28534_ (.A(_02600_),
    .B1(_02398_),
    .B2(_02924_),
    .ZN(_03348_));
 NAND2_X1 _28535_ (.A1(_02600_),
    .A2(_02602_),
    .ZN(_03349_));
 AND2_X1 _28536_ (.A1(_03348_),
    .A2(_03349_),
    .ZN(_03350_));
 OAI21_X1 _28537_ (.A(_02593_),
    .B1(_02408_),
    .B2(_02466_),
    .ZN(_03351_));
 AND4_X1 _28538_ (.A1(_03346_),
    .A2(_03347_),
    .A3(_03350_),
    .A4(_03351_),
    .ZN(_03352_));
 OAI21_X1 _28539_ (.A(_02581_),
    .B1(_02398_),
    .B2(_02404_),
    .ZN(_03353_));
 OAI21_X1 _28540_ (.A(_02575_),
    .B1(_02398_),
    .B2(_02578_),
    .ZN(_03354_));
 OAI21_X1 _28541_ (.A(_02575_),
    .B1(_02887_),
    .B2(_02455_),
    .ZN(_03355_));
 OAI21_X1 _28542_ (.A(_02581_),
    .B1(_02887_),
    .B2(_02523_),
    .ZN(_03356_));
 AND4_X1 _28543_ (.A1(_03353_),
    .A2(_03354_),
    .A3(_03355_),
    .A4(_03356_),
    .ZN(_03357_));
 AND2_X1 _28544_ (.A1(_02926_),
    .A2(_02493_),
    .ZN(_03358_));
 AND4_X1 _28545_ (.A1(_02401_),
    .A2(_02434_),
    .A3(_02417_),
    .A4(_02524_),
    .ZN(_03359_));
 OR2_X1 _28546_ (.A1(_03358_),
    .A2(_03359_),
    .ZN(_03360_));
 NAND2_X1 _28547_ (.A1(_02504_),
    .A2(_02595_),
    .ZN(_03361_));
 NAND3_X1 _28548_ (.A1(_02541_),
    .A2(_03295_),
    .A3(_02524_),
    .ZN(_03362_));
 INV_X1 _28549_ (.A(_02504_),
    .ZN(_03363_));
 OAI211_X1 _28550_ (.A(_03361_),
    .B(_03362_),
    .C1(_03308_),
    .C2(_03363_),
    .ZN(_03364_));
 AOI21_X1 _28551_ (.A(_03363_),
    .B1(_02490_),
    .B2(_02444_),
    .ZN(_03365_));
 NAND2_X1 _28552_ (.A1(_02486_),
    .A2(_02498_),
    .ZN(_03366_));
 INV_X1 _28553_ (.A(_02500_),
    .ZN(_03367_));
 INV_X1 _28554_ (.A(_02498_),
    .ZN(_03368_));
 OAI22_X1 _28555_ (.A1(_03366_),
    .A2(_02423_),
    .B1(_03367_),
    .B2(_03368_),
    .ZN(_03369_));
 NOR4_X1 _28556_ (.A1(_03360_),
    .A2(_03364_),
    .A3(_03365_),
    .A4(_03369_),
    .ZN(_03370_));
 NAND4_X1 _28557_ (.A1(_03344_),
    .A2(_03352_),
    .A3(_03357_),
    .A4(_03370_),
    .ZN(_03371_));
 NOR2_X2 _28558_ (.A1(_03338_),
    .A2(_03371_),
    .ZN(_03372_));
 OAI21_X1 _28559_ (.A(_01898_),
    .B1(_01956_),
    .B2(_01949_),
    .ZN(_03373_));
 AND2_X1 _28560_ (.A1(_01961_),
    .A2(_01903_),
    .ZN(_03374_));
 AND2_X1 _28561_ (.A1(_01960_),
    .A2(_01953_),
    .ZN(_03375_));
 AND3_X1 _28562_ (.A1(_01915_),
    .A2(_03003_),
    .A3(_01980_),
    .ZN(_03376_));
 NOR4_X1 _28563_ (.A1(_03374_),
    .A2(_02982_),
    .A3(_03375_),
    .A4(_03376_),
    .ZN(_03377_));
 OAI21_X1 _28564_ (.A(_01897_),
    .B1(_01858_),
    .B2(_02012_),
    .ZN(_03378_));
 OAI211_X1 _28565_ (.A(_01898_),
    .B(_16690_),
    .C1(_02088_),
    .C2(_01848_),
    .ZN(_03379_));
 AND4_X1 _28566_ (.A1(_03373_),
    .A2(_03377_),
    .A3(_03378_),
    .A4(_03379_),
    .ZN(_03380_));
 AND2_X1 _28567_ (.A1(_02113_),
    .A2(_01973_),
    .ZN(_03381_));
 AOI21_X1 _28568_ (.A(_03381_),
    .B1(_02971_),
    .B2(_01973_),
    .ZN(_03382_));
 NAND4_X1 _28569_ (.A1(_01852_),
    .A2(_01980_),
    .A3(_01841_),
    .A4(_01954_),
    .ZN(_03383_));
 NAND3_X1 _28570_ (.A1(_03382_),
    .A2(_02967_),
    .A3(_03383_),
    .ZN(_03384_));
 NAND2_X1 _28571_ (.A1(_02000_),
    .A2(_01983_),
    .ZN(_03385_));
 INV_X1 _28572_ (.A(_01926_),
    .ZN(_03386_));
 INV_X1 _28573_ (.A(_01949_),
    .ZN(_03387_));
 OAI211_X1 _28574_ (.A(_01930_),
    .B(_03385_),
    .C1(_03386_),
    .C2(_03387_),
    .ZN(_03388_));
 INV_X1 _28575_ (.A(_02113_),
    .ZN(_03389_));
 INV_X1 _28576_ (.A(_02037_),
    .ZN(_03390_));
 AOI21_X1 _28577_ (.A(_03386_),
    .B1(_03389_),
    .B2(_03390_),
    .ZN(_03391_));
 AND4_X1 _28578_ (.A1(_01920_),
    .A2(_01980_),
    .A3(_02061_),
    .A4(_01887_),
    .ZN(_03392_));
 NOR4_X1 _28579_ (.A1(_03384_),
    .A2(_03388_),
    .A3(_03391_),
    .A4(_03392_),
    .ZN(_03393_));
 NAND2_X1 _28580_ (.A1(_02057_),
    .A2(_01943_),
    .ZN(_03394_));
 BUF_X2 _28581_ (.A(_01943_),
    .Z(_03395_));
 OAI21_X1 _28582_ (.A(_03395_),
    .B1(_02076_),
    .B2(_01956_),
    .ZN(_03396_));
 BUF_X2 _28583_ (.A(_02018_),
    .Z(_03397_));
 OAI21_X1 _28584_ (.A(_03397_),
    .B1(_02035_),
    .B2(_02039_),
    .ZN(_03398_));
 OAI21_X1 _28585_ (.A(_03397_),
    .B1(_01947_),
    .B2(_01949_),
    .ZN(_03399_));
 AND4_X1 _28586_ (.A1(_03394_),
    .A2(_03396_),
    .A3(_03398_),
    .A4(_03399_),
    .ZN(_03400_));
 BUF_X2 _28587_ (.A(_01963_),
    .Z(_03401_));
 OAI211_X1 _28588_ (.A(_03003_),
    .B(_03020_),
    .C1(_01979_),
    .C2(_03401_),
    .ZN(_03402_));
 OAI21_X1 _28589_ (.A(_03402_),
    .B1(_02978_),
    .B2(_03023_),
    .ZN(_03403_));
 AOI211_X1 _28590_ (.A(_16690_),
    .B(_01971_),
    .C1(_02088_),
    .C2(_01848_),
    .ZN(_03404_));
 BUF_X2 _28591_ (.A(_01846_),
    .Z(_03405_));
 OAI211_X1 _28592_ (.A(_02059_),
    .B(_01905_),
    .C1(_01954_),
    .C2(_03405_),
    .ZN(_03406_));
 NAND2_X1 _28593_ (.A1(_01912_),
    .A2(_02059_),
    .ZN(_03407_));
 NAND2_X1 _28594_ (.A1(_03406_),
    .A2(_03407_),
    .ZN(_03408_));
 NAND3_X1 _28595_ (.A1(_02108_),
    .A2(_03003_),
    .A3(_03020_),
    .ZN(_03409_));
 NAND3_X1 _28596_ (.A1(_01953_),
    .A2(_02094_),
    .A3(_03020_),
    .ZN(_03410_));
 NAND3_X1 _28597_ (.A1(_03025_),
    .A2(_03409_),
    .A3(_03410_),
    .ZN(_03411_));
 NOR4_X1 _28598_ (.A1(_03403_),
    .A2(_03404_),
    .A3(_03408_),
    .A4(_03411_),
    .ZN(_03412_));
 NAND4_X1 _28599_ (.A1(_03380_),
    .A2(_03393_),
    .A3(_03400_),
    .A4(_03412_),
    .ZN(_03413_));
 AND3_X1 _28600_ (.A1(_02032_),
    .A2(_03002_),
    .A3(_01841_),
    .ZN(_03414_));
 AOI211_X1 _28601_ (.A(_02099_),
    .B(_03414_),
    .C1(_02108_),
    .C2(_01843_),
    .ZN(_03415_));
 OAI21_X1 _28602_ (.A(_01843_),
    .B1(_02971_),
    .B2(_01996_),
    .ZN(_03416_));
 OAI21_X1 _28603_ (.A(_01890_),
    .B1(_02042_),
    .B2(_02037_),
    .ZN(_03417_));
 AND4_X1 _28604_ (.A1(_01892_),
    .A2(_03415_),
    .A3(_03416_),
    .A4(_03417_),
    .ZN(_03418_));
 OAI21_X1 _28605_ (.A(_02047_),
    .B1(_02032_),
    .B2(_02033_),
    .ZN(_03419_));
 OAI21_X1 _28606_ (.A(_02014_),
    .B1(_02032_),
    .B2(_01858_),
    .ZN(_03420_));
 OAI21_X1 _28607_ (.A(_02014_),
    .B1(_02113_),
    .B2(_02039_),
    .ZN(_03421_));
 OAI21_X1 _28608_ (.A(_02047_),
    .B1(_02113_),
    .B2(_03401_),
    .ZN(_03422_));
 AND4_X1 _28609_ (.A1(_03419_),
    .A2(_03420_),
    .A3(_03421_),
    .A4(_03422_),
    .ZN(_03423_));
 MUX2_X1 _28610_ (.A(_01938_),
    .B(_01867_),
    .S(_01881_),
    .Z(_03424_));
 AND2_X1 _28611_ (.A1(_03424_),
    .A2(_01958_),
    .ZN(_03425_));
 INV_X1 _28612_ (.A(_02000_),
    .ZN(_03426_));
 AOI21_X1 _28613_ (.A(_02125_),
    .B1(_03426_),
    .B2(_01944_),
    .ZN(_03427_));
 NAND3_X1 _28614_ (.A1(_01915_),
    .A2(_03003_),
    .A3(_01932_),
    .ZN(_03428_));
 NAND3_X1 _28615_ (.A1(_02129_),
    .A2(_02127_),
    .A3(_03428_),
    .ZN(_03429_));
 NAND2_X1 _28616_ (.A1(_02007_),
    .A2(_01957_),
    .ZN(_03430_));
 INV_X1 _28617_ (.A(_01992_),
    .ZN(_03431_));
 OAI22_X1 _28618_ (.A1(_03430_),
    .A2(_01856_),
    .B1(_02068_),
    .B2(_03431_),
    .ZN(_03432_));
 NOR4_X1 _28619_ (.A1(_03425_),
    .A2(_03427_),
    .A3(_03429_),
    .A4(_03432_),
    .ZN(_03433_));
 OAI21_X1 _28620_ (.A(_02132_),
    .B1(_02001_),
    .B2(_02039_),
    .ZN(_03434_));
 NAND4_X1 _28621_ (.A1(_01887_),
    .A2(_02103_),
    .A3(_01932_),
    .A4(_02088_),
    .ZN(_03435_));
 NAND3_X1 _28622_ (.A1(_02132_),
    .A2(_01935_),
    .A3(_02009_),
    .ZN(_03436_));
 NAND3_X1 _28623_ (.A1(_03434_),
    .A2(_03435_),
    .A3(_03436_),
    .ZN(_03437_));
 NAND2_X1 _28624_ (.A1(_01934_),
    .A2(_02037_),
    .ZN(_03438_));
 INV_X1 _28625_ (.A(_01933_),
    .ZN(_03439_));
 OAI211_X1 _28626_ (.A(_03438_),
    .B(_01967_),
    .C1(_03389_),
    .C2(_03439_),
    .ZN(_03440_));
 AOI21_X1 _28627_ (.A(_03439_),
    .B1(_02068_),
    .B2(_03387_),
    .ZN(_03441_));
 NOR2_X1 _28628_ (.A1(_01927_),
    .A2(_01894_),
    .ZN(_03442_));
 AND2_X1 _28629_ (.A1(_01934_),
    .A2(_03442_),
    .ZN(_03443_));
 NOR4_X1 _28630_ (.A1(_03437_),
    .A2(_03440_),
    .A3(_03441_),
    .A4(_03443_),
    .ZN(_03444_));
 NAND4_X1 _28631_ (.A1(_03418_),
    .A2(_03423_),
    .A3(_03433_),
    .A4(_03444_),
    .ZN(_03445_));
 NOR2_X2 _28632_ (.A1(_03413_),
    .A2(_03445_),
    .ZN(_03446_));
 XNOR2_X1 _28633_ (.A(_03372_),
    .B(_03446_),
    .ZN(_03447_));
 NAND2_X1 _28634_ (.A1(_02330_),
    .A2(_02361_),
    .ZN(_03448_));
 AND3_X1 _28635_ (.A1(_02194_),
    .A2(_02260_),
    .A3(_02227_),
    .ZN(_03449_));
 AOI211_X1 _28636_ (.A(_03449_),
    .B(_03066_),
    .C1(_02223_),
    .C2(_02334_),
    .ZN(_03450_));
 OAI21_X1 _28637_ (.A(_02152_),
    .B1(_02214_),
    .B2(_02353_),
    .ZN(_03451_));
 OAI211_X1 _28638_ (.A(_02152_),
    .B(_16770_),
    .C1(_02375_),
    .C2(_02182_),
    .ZN(_03452_));
 AND4_X1 _28639_ (.A1(_03448_),
    .A2(_03450_),
    .A3(_03451_),
    .A4(_03452_),
    .ZN(_03453_));
 NOR2_X1 _28640_ (.A1(_02143_),
    .A2(_02188_),
    .ZN(_03454_));
 AND2_X1 _28641_ (.A1(_03454_),
    .A2(_02234_),
    .ZN(_03455_));
 INV_X1 _28642_ (.A(_03455_),
    .ZN(_03456_));
 NAND3_X1 _28643_ (.A1(_02235_),
    .A2(_02174_),
    .A3(_03061_),
    .ZN(_03457_));
 INV_X1 _28644_ (.A(_02368_),
    .ZN(_03458_));
 INV_X1 _28645_ (.A(_02234_),
    .ZN(_03459_));
 OAI211_X1 _28646_ (.A(_03456_),
    .B(_03457_),
    .C1(_03458_),
    .C2(_03459_),
    .ZN(_03460_));
 INV_X1 _28647_ (.A(_02274_),
    .ZN(_03461_));
 INV_X1 _28648_ (.A(_02378_),
    .ZN(_03462_));
 INV_X1 _28649_ (.A(_02276_),
    .ZN(_03463_));
 AOI21_X1 _28650_ (.A(_03461_),
    .B1(_03462_),
    .B2(_03463_),
    .ZN(_03464_));
 AND3_X1 _28651_ (.A1(_02278_),
    .A2(_02308_),
    .A3(_02239_),
    .ZN(_03465_));
 NOR4_X1 _28652_ (.A1(_03460_),
    .A2(_03126_),
    .A3(_03464_),
    .A4(_03465_),
    .ZN(_03466_));
 NAND2_X1 _28653_ (.A1(_03062_),
    .A2(_02245_),
    .ZN(_03467_));
 NAND3_X1 _28654_ (.A1(_02368_),
    .A2(_02260_),
    .A3(_02261_),
    .ZN(_03468_));
 OAI21_X1 _28655_ (.A(_02245_),
    .B1(_03056_),
    .B2(_02361_),
    .ZN(_03469_));
 OAI211_X1 _28656_ (.A(_02260_),
    .B(_02261_),
    .C1(_02356_),
    .C2(_02333_),
    .ZN(_03470_));
 NAND4_X1 _28657_ (.A1(_03467_),
    .A2(_03468_),
    .A3(_03469_),
    .A4(_03470_),
    .ZN(_03471_));
 NAND2_X1 _28658_ (.A1(_02200_),
    .A2(_02265_),
    .ZN(_03472_));
 NAND3_X1 _28659_ (.A1(_02265_),
    .A2(_02352_),
    .A3(_02174_),
    .ZN(_03473_));
 NAND2_X1 _28660_ (.A1(_03472_),
    .A2(_03473_),
    .ZN(_03474_));
 NAND2_X1 _28661_ (.A1(_02311_),
    .A2(_02263_),
    .ZN(_03475_));
 NAND3_X1 _28662_ (.A1(_02265_),
    .A2(_02198_),
    .A3(_02353_),
    .ZN(_03476_));
 NAND3_X1 _28663_ (.A1(_02265_),
    .A2(_03075_),
    .A3(_02353_),
    .ZN(_03477_));
 NAND3_X1 _28664_ (.A1(_03475_),
    .A2(_03476_),
    .A3(_03477_),
    .ZN(_03478_));
 NOR4_X1 _28665_ (.A1(_03471_),
    .A2(_02302_),
    .A3(_03474_),
    .A4(_03478_),
    .ZN(_03479_));
 OAI211_X1 _28666_ (.A(_03052_),
    .B(_02353_),
    .C1(_02375_),
    .C2(_03080_),
    .ZN(_03480_));
 OAI211_X1 _28667_ (.A(_03052_),
    .B(_02352_),
    .C1(_02375_),
    .C2(_03080_),
    .ZN(_03481_));
 OAI21_X1 _28668_ (.A(_03052_),
    .B1(_02288_),
    .B2(_02356_),
    .ZN(_03482_));
 OAI21_X1 _28669_ (.A(_03052_),
    .B1(_02347_),
    .B2(_02361_),
    .ZN(_03483_));
 NAND4_X1 _28670_ (.A1(_03480_),
    .A2(_03481_),
    .A3(_03482_),
    .A4(_03483_),
    .ZN(_03484_));
 INV_X1 _28671_ (.A(_02219_),
    .ZN(_03485_));
 OAI21_X1 _28672_ (.A(_03055_),
    .B1(_03485_),
    .B2(_03458_),
    .ZN(_03486_));
 AND2_X1 _28673_ (.A1(_02254_),
    .A2(_02219_),
    .ZN(_03487_));
 AND3_X1 _28674_ (.A1(_02146_),
    .A2(_02220_),
    .A3(_02259_),
    .ZN(_03488_));
 NOR4_X1 _28675_ (.A1(_03484_),
    .A2(_03486_),
    .A3(_03487_),
    .A4(_03488_),
    .ZN(_03489_));
 NAND4_X1 _28676_ (.A1(_03453_),
    .A2(_03466_),
    .A3(_03479_),
    .A4(_03489_),
    .ZN(_03490_));
 INV_X1 _28677_ (.A(_02322_),
    .ZN(_03491_));
 INV_X1 _28678_ (.A(_02215_),
    .ZN(_03492_));
 OAI211_X1 _28679_ (.A(_03491_),
    .B(_02346_),
    .C1(_03072_),
    .C2(_03492_),
    .ZN(_03493_));
 NAND2_X1 _28680_ (.A1(_02215_),
    .A2(_02200_),
    .ZN(_03494_));
 NAND2_X1 _28681_ (.A1(_02343_),
    .A2(_03494_),
    .ZN(_03495_));
 OAI21_X1 _28682_ (.A(_02192_),
    .B1(_02336_),
    .B2(_02318_),
    .ZN(_03496_));
 NAND2_X1 _28683_ (.A1(_02191_),
    .A2(_02199_),
    .ZN(_03497_));
 OAI211_X1 _28684_ (.A(_03496_),
    .B(_03497_),
    .C1(_03114_),
    .C2(_02250_),
    .ZN(_03498_));
 NOR4_X1 _28685_ (.A1(_03493_),
    .A2(_03495_),
    .A3(_02210_),
    .A4(_03498_),
    .ZN(_03499_));
 NOR2_X1 _28686_ (.A1(_02248_),
    .A2(_03056_),
    .ZN(_03500_));
 AOI21_X1 _28687_ (.A(_02376_),
    .B1(_03500_),
    .B2(_03458_),
    .ZN(_03501_));
 NAND2_X1 _28688_ (.A1(_03454_),
    .A2(_02380_),
    .ZN(_03502_));
 NAND3_X1 _28689_ (.A1(_02380_),
    .A2(_02352_),
    .A3(_02188_),
    .ZN(_03503_));
 NAND2_X1 _28690_ (.A1(_03502_),
    .A2(_03503_),
    .ZN(_03504_));
 NOR2_X1 _28691_ (.A1(_03501_),
    .A2(_03504_),
    .ZN(_03505_));
 OAI21_X1 _28692_ (.A(_02326_),
    .B1(_02363_),
    .B2(_02318_),
    .ZN(_03506_));
 NAND3_X1 _28693_ (.A1(_02222_),
    .A2(_02179_),
    .A3(_02171_),
    .ZN(_03507_));
 OAI211_X1 _28694_ (.A(_02326_),
    .B(_02352_),
    .C1(_02375_),
    .C2(_02285_),
    .ZN(_03508_));
 AND4_X1 _28695_ (.A1(_03505_),
    .A2(_03506_),
    .A3(_03507_),
    .A4(_03508_),
    .ZN(_03509_));
 OAI21_X1 _28696_ (.A(_02369_),
    .B1(_02246_),
    .B2(_02248_),
    .ZN(_03510_));
 OAI21_X1 _28697_ (.A(_02212_),
    .B1(_02246_),
    .B2(_02318_),
    .ZN(_03511_));
 OAI21_X1 _28698_ (.A(_02212_),
    .B1(_02254_),
    .B2(_02276_),
    .ZN(_03512_));
 OAI21_X1 _28699_ (.A(_02369_),
    .B1(_02254_),
    .B2(_02333_),
    .ZN(_03513_));
 AND4_X1 _28700_ (.A1(_03510_),
    .A2(_03511_),
    .A3(_03512_),
    .A4(_03513_),
    .ZN(_03514_));
 OAI21_X1 _28701_ (.A(_02339_),
    .B1(_03061_),
    .B2(_02221_),
    .ZN(_03515_));
 NAND2_X1 _28702_ (.A1(_02339_),
    .A2(_02268_),
    .ZN(_03516_));
 NAND2_X1 _28703_ (.A1(_02292_),
    .A2(_02368_),
    .ZN(_03517_));
 NAND2_X1 _28704_ (.A1(_02339_),
    .A2(_02214_),
    .ZN(_03518_));
 AND3_X1 _28705_ (.A1(_03516_),
    .A2(_03517_),
    .A3(_03518_),
    .ZN(_03519_));
 OAI21_X1 _28706_ (.A(_02358_),
    .B1(_02328_),
    .B2(_02370_),
    .ZN(_03520_));
 OAI21_X1 _28707_ (.A(_02358_),
    .B1(_02204_),
    .B2(_02276_),
    .ZN(_03521_));
 AND4_X1 _28708_ (.A1(_03515_),
    .A2(_03519_),
    .A3(_03520_),
    .A4(_03521_),
    .ZN(_03522_));
 NAND4_X1 _28709_ (.A1(_03499_),
    .A2(_03509_),
    .A3(_03514_),
    .A4(_03522_),
    .ZN(_03523_));
 NOR2_X2 _28710_ (.A1(_03490_),
    .A2(_03523_),
    .ZN(_03524_));
 XNOR2_X1 _28711_ (.A(_03447_),
    .B(_03524_),
    .ZN(_03525_));
 NAND3_X1 _28712_ (.A1(_03175_),
    .A2(_02638_),
    .A3(_03246_),
    .ZN(_03526_));
 NAND3_X1 _28713_ (.A1(_03175_),
    .A2(_02684_),
    .A3(_03246_),
    .ZN(_03527_));
 BUF_X2 _28714_ (.A(_02627_),
    .Z(_03528_));
 NAND3_X1 _28715_ (.A1(_03175_),
    .A2(_03528_),
    .A3(_03246_),
    .ZN(_03529_));
 NAND3_X1 _28716_ (.A1(_03526_),
    .A2(_03527_),
    .A3(_03529_),
    .ZN(_03530_));
 AND2_X1 _28717_ (.A1(_02727_),
    .A2(_03175_),
    .ZN(_03531_));
 AND2_X1 _28718_ (.A1(_02679_),
    .A2(_02674_),
    .ZN(_03532_));
 AND2_X1 _28719_ (.A1(_02680_),
    .A2(_03156_),
    .ZN(_03533_));
 NOR4_X1 _28720_ (.A1(_03530_),
    .A2(_03531_),
    .A3(_03532_),
    .A4(_03533_),
    .ZN(_03534_));
 INV_X1 _28721_ (.A(_02736_),
    .ZN(_03535_));
 NAND2_X1 _28722_ (.A1(_02761_),
    .A2(_02748_),
    .ZN(_03536_));
 NOR2_X1 _28723_ (.A1(_03535_),
    .A2(_03536_),
    .ZN(_03537_));
 NAND2_X1 _28724_ (.A1(_02742_),
    .A2(_02815_),
    .ZN(_03538_));
 NAND2_X1 _28725_ (.A1(_02739_),
    .A2(_03538_),
    .ZN(_03539_));
 AOI211_X1 _28726_ (.A(_03537_),
    .B(_03539_),
    .C1(_02793_),
    .C2(_02742_),
    .ZN(_03540_));
 BUF_X2 _28727_ (.A(_02695_),
    .Z(_03541_));
 NAND2_X1 _28728_ (.A1(_03541_),
    .A2(_02727_),
    .ZN(_03542_));
 NAND2_X1 _28729_ (.A1(_02682_),
    .A2(_02695_),
    .ZN(_03543_));
 AND2_X1 _28730_ (.A1(_02748_),
    .A2(_02829_),
    .ZN(_03544_));
 NAND2_X1 _28731_ (.A1(_03541_),
    .A2(_03544_),
    .ZN(_03545_));
 AND4_X1 _28732_ (.A1(_03542_),
    .A2(_03543_),
    .A3(_03545_),
    .A4(_02697_),
    .ZN(_03546_));
 NAND3_X1 _28733_ (.A1(_02733_),
    .A2(_02800_),
    .A3(_03528_),
    .ZN(_03547_));
 OAI21_X1 _28734_ (.A(_02733_),
    .B1(_03169_),
    .B2(_03209_),
    .ZN(_03548_));
 BUF_X2 _28735_ (.A(_02702_),
    .Z(_03549_));
 OAI211_X1 _28736_ (.A(_02733_),
    .B(_03549_),
    .C1(_02747_),
    .C2(_02657_),
    .ZN(_03550_));
 AND4_X1 _28737_ (.A1(_03547_),
    .A2(_03144_),
    .A3(_03548_),
    .A4(_03550_),
    .ZN(_03551_));
 AND4_X1 _28738_ (.A1(_03534_),
    .A2(_03540_),
    .A3(_03546_),
    .A4(_03551_),
    .ZN(_03552_));
 OAI21_X1 _28739_ (.A(_03204_),
    .B1(_02818_),
    .B2(_03209_),
    .ZN(_03553_));
 NAND2_X1 _28740_ (.A1(_02765_),
    .A2(_03204_),
    .ZN(_03554_));
 AND2_X1 _28741_ (.A1(_02796_),
    .A2(_03204_),
    .ZN(_03555_));
 INV_X1 _28742_ (.A(_03555_),
    .ZN(_03556_));
 AND4_X1 _28743_ (.A1(_02791_),
    .A2(_03553_),
    .A3(_03554_),
    .A4(_03556_),
    .ZN(_03557_));
 CLKBUF_X2 _28744_ (.A(_02630_),
    .Z(_03558_));
 AND2_X1 _28745_ (.A1(_03558_),
    .A2(_02780_),
    .ZN(_03559_));
 AOI211_X1 _28746_ (.A(_16778_),
    .B(_03206_),
    .C1(_02829_),
    .C2(_02650_),
    .ZN(_03560_));
 AOI221_X4 _28747_ (.A(_03559_),
    .B1(_02780_),
    .B2(_02809_),
    .C1(_03560_),
    .C2(_02743_),
    .ZN(_03561_));
 AND2_X1 _28748_ (.A1(_03558_),
    .A2(_03172_),
    .ZN(_03562_));
 AND2_X1 _28749_ (.A1(_02782_),
    .A2(_02769_),
    .ZN(_03563_));
 AND2_X1 _28750_ (.A1(_02769_),
    .A2(_02813_),
    .ZN(_03564_));
 NOR4_X1 _28751_ (.A1(_02768_),
    .A2(_03562_),
    .A3(_03563_),
    .A4(_03564_),
    .ZN(_03565_));
 OAI21_X1 _28752_ (.A(_02759_),
    .B1(_02796_),
    .B2(_02671_),
    .ZN(_03566_));
 NAND3_X1 _28753_ (.A1(_02759_),
    .A2(_02638_),
    .A3(_02748_),
    .ZN(_03567_));
 NAND2_X1 _28754_ (.A1(_02782_),
    .A2(_02759_),
    .ZN(_03568_));
 AND4_X1 _28755_ (.A1(_03177_),
    .A2(_03566_),
    .A3(_03567_),
    .A4(_03568_),
    .ZN(_03569_));
 AND4_X1 _28756_ (.A1(_03557_),
    .A2(_03561_),
    .A3(_03565_),
    .A4(_03569_),
    .ZN(_03570_));
 INV_X1 _28757_ (.A(_02641_),
    .ZN(_03571_));
 INV_X1 _28758_ (.A(_02682_),
    .ZN(_03572_));
 AOI21_X1 _28759_ (.A(_03146_),
    .B1(_03571_),
    .B2(_03572_),
    .ZN(_03573_));
 INV_X1 _28760_ (.A(_03536_),
    .ZN(_03574_));
 NAND2_X1 _28761_ (.A1(_03574_),
    .A2(_02723_),
    .ZN(_03575_));
 INV_X1 _28762_ (.A(_03575_),
    .ZN(_03576_));
 AND2_X1 _28763_ (.A1(_02723_),
    .A2(_03549_),
    .ZN(_03577_));
 AND4_X1 _28764_ (.A1(_02747_),
    .A2(_02622_),
    .A3(_02676_),
    .A4(_02667_),
    .ZN(_03578_));
 NOR4_X1 _28765_ (.A1(_03573_),
    .A2(_03576_),
    .A3(_03577_),
    .A4(_03578_),
    .ZN(_03579_));
 AND2_X1 _28766_ (.A1(_03169_),
    .A2(_02664_),
    .ZN(_03580_));
 INV_X1 _28767_ (.A(_02664_),
    .ZN(_03581_));
 AOI21_X1 _28768_ (.A(_03581_),
    .B1(_03152_),
    .B2(_03572_),
    .ZN(_03582_));
 AOI211_X1 _28769_ (.A(_03580_),
    .B(_03582_),
    .C1(_02665_),
    .C2(_03544_),
    .ZN(_03583_));
 AOI21_X1 _28770_ (.A(_02713_),
    .B1(_02817_),
    .B2(_02688_),
    .ZN(_03584_));
 AOI21_X1 _28771_ (.A(_02713_),
    .B1(_02807_),
    .B2(_02808_),
    .ZN(_03585_));
 AND2_X1 _28772_ (.A1(_02709_),
    .A2(_02813_),
    .ZN(_03586_));
 AND2_X1 _28773_ (.A1(_02709_),
    .A2(_03558_),
    .ZN(_03587_));
 NOR4_X1 _28774_ (.A1(_03584_),
    .A2(_03585_),
    .A3(_03586_),
    .A4(_03587_),
    .ZN(_03588_));
 NAND4_X1 _28775_ (.A1(_02622_),
    .A2(_02684_),
    .A3(_03246_),
    .A4(_03234_),
    .ZN(_03589_));
 OAI21_X1 _28776_ (.A(_02635_),
    .B1(_03558_),
    .B2(_02670_),
    .ZN(_03590_));
 AND4_X1 _28777_ (.A1(_02649_),
    .A2(_02644_),
    .A3(_03589_),
    .A4(_03590_),
    .ZN(_03591_));
 AND4_X1 _28778_ (.A1(_03579_),
    .A2(_03583_),
    .A3(_03588_),
    .A4(_03591_),
    .ZN(_03592_));
 NAND2_X1 _28779_ (.A1(_02828_),
    .A2(_02813_),
    .ZN(_03593_));
 AND2_X1 _28780_ (.A1(_02821_),
    .A2(_02796_),
    .ZN(_03594_));
 INV_X1 _28781_ (.A(_03594_),
    .ZN(_03595_));
 NAND2_X1 _28782_ (.A1(_02711_),
    .A2(_02828_),
    .ZN(_03596_));
 OAI21_X1 _28783_ (.A(_02828_),
    .B1(_02724_),
    .B2(_03156_),
    .ZN(_03597_));
 AND4_X1 _28784_ (.A1(_03593_),
    .A2(_03595_),
    .A3(_03596_),
    .A4(_03597_),
    .ZN(_03598_));
 NAND3_X1 _28785_ (.A1(_03237_),
    .A2(_03211_),
    .A3(_03234_),
    .ZN(_03599_));
 OAI21_X1 _28786_ (.A(_02831_),
    .B1(_03150_),
    .B2(_03203_),
    .ZN(_03600_));
 NAND2_X1 _28787_ (.A1(_02782_),
    .A2(_02831_),
    .ZN(_03601_));
 NAND4_X1 _28788_ (.A1(_03598_),
    .A2(_03599_),
    .A3(_03600_),
    .A4(_03601_),
    .ZN(_03602_));
 INV_X1 _28789_ (.A(_02812_),
    .ZN(_03603_));
 AOI21_X1 _28790_ (.A(_03603_),
    .B1(_02719_),
    .B2(_02807_),
    .ZN(_03604_));
 AND2_X1 _28791_ (.A1(_02805_),
    .A2(_02658_),
    .ZN(_03605_));
 AND2_X1 _28792_ (.A1(_02805_),
    .A2(_02698_),
    .ZN(_03606_));
 AND2_X1 _28793_ (.A1(_02805_),
    .A2(_02800_),
    .ZN(_03607_));
 AND2_X1 _28794_ (.A1(_02804_),
    .A2(_02632_),
    .ZN(_03608_));
 OR4_X1 _28795_ (.A1(_03605_),
    .A2(_03606_),
    .A3(_03607_),
    .A4(_03608_),
    .ZN(_03609_));
 NAND4_X1 _28796_ (.A1(_03211_),
    .A2(_03528_),
    .A3(_02676_),
    .A4(_02667_),
    .ZN(_03610_));
 NAND2_X1 _28797_ (.A1(_03243_),
    .A2(_03610_),
    .ZN(_03611_));
 NOR4_X1 _28798_ (.A1(_03602_),
    .A2(_03604_),
    .A3(_03609_),
    .A4(_03611_),
    .ZN(_03612_));
 AND4_X1 _28799_ (.A1(_03552_),
    .A2(_03570_),
    .A3(_03592_),
    .A4(_03612_),
    .ZN(_03613_));
 INV_X1 _28800_ (.A(_03199_),
    .ZN(_03614_));
 NAND2_X2 _28801_ (.A1(_03613_),
    .A2(_03614_),
    .ZN(_03615_));
 XNOR2_X1 _28802_ (.A(_03615_),
    .B(_03042_),
    .ZN(_03616_));
 XNOR2_X1 _28803_ (.A(_03525_),
    .B(_03616_),
    .ZN(_03617_));
 INV_X1 _28804_ (.A(_17153_),
    .ZN(_03618_));
 XNOR2_X1 _28805_ (.A(_03617_),
    .B(_03618_),
    .ZN(_03619_));
 MUX2_X1 _28806_ (.A(_03290_),
    .B(_03619_),
    .S(_01825_),
    .Z(_00710_));
 XOR2_X1 _28807_ (.A(_17113_),
    .B(_17177_),
    .Z(_03620_));
 XOR2_X1 _28808_ (.A(_17081_),
    .B(_17145_),
    .Z(_03621_));
 XNOR2_X1 _28809_ (.A(_03620_),
    .B(_03621_),
    .ZN(_03622_));
 XOR2_X1 _28810_ (.A(_16110_),
    .B(_03622_),
    .Z(_03623_));
 MUX2_X1 _28811_ (.A(_01244_),
    .B(_03623_),
    .S(_03265_),
    .Z(_01168_));
 XOR2_X1 _28812_ (.A(_17114_),
    .B(_17178_),
    .Z(_03624_));
 XOR2_X1 _28813_ (.A(_17082_),
    .B(_17146_),
    .Z(_03625_));
 XNOR2_X1 _28814_ (.A(_03624_),
    .B(_03625_),
    .ZN(_03626_));
 XOR2_X1 _28815_ (.A(_16160_),
    .B(_03626_),
    .Z(_03627_));
 MUX2_X1 _28816_ (.A(_01245_),
    .B(_03627_),
    .S(_03265_),
    .Z(_01169_));
 XNOR2_X1 _28817_ (.A(_11040_),
    .B(_01013_),
    .ZN(_03628_));
 XNOR2_X1 _28818_ (.A(_03628_),
    .B(_17115_),
    .ZN(_03629_));
 XOR2_X1 _28819_ (.A(_17147_),
    .B(_17179_),
    .Z(_03630_));
 XOR2_X1 _28820_ (.A(_03629_),
    .B(_03630_),
    .Z(_03631_));
 XNOR2_X1 _28821_ (.A(_16408_),
    .B(_03631_),
    .ZN(_03632_));
 MUX2_X1 _28822_ (.A(_01246_),
    .B(_03632_),
    .S(_01736_),
    .Z(_01170_));
 XNOR2_X1 _28823_ (.A(_11046_),
    .B(_01015_),
    .ZN(_03633_));
 XNOR2_X1 _28824_ (.A(_03633_),
    .B(_17116_),
    .ZN(_03634_));
 XNOR2_X1 _28825_ (.A(_17148_),
    .B(_17180_),
    .ZN(_03635_));
 XOR2_X1 _28826_ (.A(_03634_),
    .B(_03635_),
    .Z(_03636_));
 XNOR2_X1 _28827_ (.A(_16518_),
    .B(_03636_),
    .ZN(_03637_));
 MUX2_X1 _28828_ (.A(_01247_),
    .B(_03637_),
    .S(_01736_),
    .Z(_01171_));
 XNOR2_X1 _28829_ (.A(_17085_),
    .B(_01017_),
    .ZN(_03638_));
 INV_X1 _28830_ (.A(_17117_),
    .ZN(_03639_));
 XNOR2_X1 _28831_ (.A(_03638_),
    .B(_03639_),
    .ZN(_03640_));
 XOR2_X1 _28832_ (.A(_17149_),
    .B(_17181_),
    .Z(_03641_));
 XOR2_X1 _28833_ (.A(_03640_),
    .B(_03641_),
    .Z(_03642_));
 XNOR2_X1 _28834_ (.A(_16608_),
    .B(_03642_),
    .ZN(_03643_));
 MUX2_X1 _28835_ (.A(_01248_),
    .B(_03643_),
    .S(_01736_),
    .Z(_01172_));
 XNOR2_X1 _28836_ (.A(_17086_),
    .B(_01019_),
    .ZN(_03644_));
 XNOR2_X1 _28837_ (.A(_03644_),
    .B(_17118_),
    .ZN(_03645_));
 XOR2_X1 _28838_ (.A(_17150_),
    .B(_17182_),
    .Z(_03646_));
 XNOR2_X1 _28839_ (.A(_03645_),
    .B(_03646_),
    .ZN(_03647_));
 XNOR2_X1 _28840_ (.A(_01341_),
    .B(_03647_),
    .ZN(_03648_));
 MUX2_X1 _28841_ (.A(_01249_),
    .B(_03648_),
    .S(_01736_),
    .Z(_01173_));
 XNOR2_X1 _28842_ (.A(_17087_),
    .B(_01021_),
    .ZN(_03649_));
 XNOR2_X1 _28843_ (.A(_03649_),
    .B(_17119_),
    .ZN(_03650_));
 XNOR2_X1 _28844_ (.A(_17151_),
    .B(_17183_),
    .ZN(_03651_));
 XOR2_X1 _28845_ (.A(_03650_),
    .B(_03651_),
    .Z(_03652_));
 XNOR2_X1 _28846_ (.A(_01404_),
    .B(_03652_),
    .ZN(_03653_));
 MUX2_X1 _28847_ (.A(_01250_),
    .B(_03653_),
    .S(_01736_),
    .Z(_01174_));
 XOR2_X1 _28848_ (.A(_17088_),
    .B(_01023_),
    .Z(_03654_));
 XNOR2_X1 _28849_ (.A(_03654_),
    .B(_17120_),
    .ZN(_03655_));
 XOR2_X1 _28850_ (.A(_17152_),
    .B(_17184_),
    .Z(_03656_));
 XOR2_X1 _28851_ (.A(_03655_),
    .B(_03656_),
    .Z(_03657_));
 XNOR2_X1 _28852_ (.A(_01466_),
    .B(_03657_),
    .ZN(_03658_));
 MUX2_X1 _28853_ (.A(_01251_),
    .B(_03658_),
    .S(_01736_),
    .Z(_01175_));
 XNOR2_X1 _28854_ (.A(_17090_),
    .B(_01025_),
    .ZN(_03659_));
 XNOR2_X1 _28855_ (.A(_03659_),
    .B(_17122_),
    .ZN(_03660_));
 XOR2_X1 _28856_ (.A(_17154_),
    .B(_17186_),
    .Z(_03661_));
 XNOR2_X1 _28857_ (.A(_03660_),
    .B(_03661_),
    .ZN(_03662_));
 XNOR2_X1 _28858_ (.A(_01517_),
    .B(_03662_),
    .ZN(_03663_));
 MUX2_X1 _28859_ (.A(_01253_),
    .B(_03663_),
    .S(_01736_),
    .Z(_01177_));
 XOR2_X1 _28860_ (.A(_17091_),
    .B(_01027_),
    .Z(_03664_));
 XNOR2_X1 _28861_ (.A(_03664_),
    .B(_17123_),
    .ZN(_03665_));
 XOR2_X1 _28862_ (.A(_17155_),
    .B(_17187_),
    .Z(_03666_));
 XOR2_X1 _28863_ (.A(_03665_),
    .B(_03666_),
    .Z(_03667_));
 XNOR2_X1 _28864_ (.A(_01567_),
    .B(_03667_),
    .ZN(_03668_));
 MUX2_X1 _28865_ (.A(_01254_),
    .B(_03668_),
    .S(_01736_),
    .Z(_01178_));
 XOR2_X1 _28866_ (.A(_17156_),
    .B(_17026_),
    .Z(_03669_));
 XOR2_X2 _28867_ (.A(_02139_),
    .B(_03446_),
    .Z(_03670_));
 NAND4_X1 _28868_ (.A1(_02227_),
    .A2(_02285_),
    .A3(_02178_),
    .A4(_02162_),
    .ZN(_03671_));
 NAND2_X1 _28869_ (.A1(_02219_),
    .A2(_02167_),
    .ZN(_03672_));
 AND2_X1 _28870_ (.A1(_02219_),
    .A2(_02311_),
    .ZN(_03673_));
 AND2_X1 _28871_ (.A1(_02219_),
    .A2(_02344_),
    .ZN(_03674_));
 NOR2_X1 _28872_ (.A1(_03673_),
    .A2(_03674_),
    .ZN(_03675_));
 INV_X1 _28873_ (.A(_03487_),
    .ZN(_03676_));
 AND4_X1 _28874_ (.A1(_03672_),
    .A2(_03675_),
    .A3(_03058_),
    .A4(_03676_),
    .ZN(_03677_));
 OAI211_X1 _28875_ (.A(_02238_),
    .B(_02240_),
    .C1(_03075_),
    .C2(_03080_),
    .ZN(_03678_));
 AND4_X1 _28876_ (.A1(_02271_),
    .A2(_02148_),
    .A3(_02178_),
    .A4(_02275_),
    .ZN(_03679_));
 AOI211_X1 _28877_ (.A(_03679_),
    .B(_03051_),
    .C1(_02206_),
    .C2(_02238_),
    .ZN(_03680_));
 AND4_X1 _28878_ (.A1(_03671_),
    .A2(_03677_),
    .A3(_03678_),
    .A4(_03680_),
    .ZN(_03681_));
 OAI211_X1 _28879_ (.A(_02308_),
    .B(_02225_),
    .C1(_02271_),
    .C2(_02285_),
    .ZN(_03682_));
 OAI211_X1 _28880_ (.A(_02308_),
    .B(_02240_),
    .C1(_02166_),
    .C2(_02145_),
    .ZN(_03683_));
 OAI21_X1 _28881_ (.A(_02308_),
    .B1(_02347_),
    .B2(_02361_),
    .ZN(_03684_));
 NAND2_X1 _28882_ (.A1(_02288_),
    .A2(_02308_),
    .ZN(_03685_));
 NAND4_X1 _28883_ (.A1(_03682_),
    .A2(_03683_),
    .A3(_03684_),
    .A4(_03685_),
    .ZN(_03686_));
 OAI211_X1 _28884_ (.A(_02234_),
    .B(_02162_),
    .C1(_02198_),
    .C2(_02188_),
    .ZN(_03687_));
 NAND3_X1 _28885_ (.A1(_03687_),
    .A2(_02269_),
    .A3(_03133_),
    .ZN(_03688_));
 INV_X1 _28886_ (.A(_02332_),
    .ZN(_03689_));
 AOI21_X1 _28887_ (.A(_03459_),
    .B1(_02357_),
    .B2(_03689_),
    .ZN(_03690_));
 NAND2_X1 _28888_ (.A1(_02194_),
    .A2(_02234_),
    .ZN(_03691_));
 OAI21_X1 _28889_ (.A(_03691_),
    .B1(_03459_),
    .B2(_02250_),
    .ZN(_03692_));
 NOR4_X1 _28890_ (.A1(_03686_),
    .A2(_03688_),
    .A3(_03690_),
    .A4(_03692_),
    .ZN(_03693_));
 OAI21_X1 _28891_ (.A(_02263_),
    .B1(_02222_),
    .B2(_02332_),
    .ZN(_03694_));
 OAI211_X1 _28892_ (.A(_02263_),
    .B(_02157_),
    .C1(_02375_),
    .C2(_02158_),
    .ZN(_03695_));
 OAI21_X1 _28893_ (.A(_02263_),
    .B1(_02317_),
    .B2(_02294_),
    .ZN(_03696_));
 AND4_X1 _28894_ (.A1(_03475_),
    .A2(_03694_),
    .A3(_03695_),
    .A4(_03696_),
    .ZN(_03697_));
 NAND2_X1 _28895_ (.A1(_02245_),
    .A2(_02333_),
    .ZN(_03698_));
 OR2_X1 _28896_ (.A1(_02344_),
    .A2(_02311_),
    .ZN(_03699_));
 OAI21_X1 _28897_ (.A(_02245_),
    .B1(_03699_),
    .B2(_03056_),
    .ZN(_03700_));
 AND4_X1 _28898_ (.A1(_02256_),
    .A2(_03697_),
    .A3(_03698_),
    .A4(_03700_),
    .ZN(_03701_));
 OAI21_X1 _28899_ (.A(_02152_),
    .B1(_02311_),
    .B2(_02214_),
    .ZN(_03702_));
 AND2_X1 _28900_ (.A1(_02146_),
    .A2(_02259_),
    .ZN(_03703_));
 OAI21_X1 _28901_ (.A(_02151_),
    .B1(_03703_),
    .B2(_02379_),
    .ZN(_03704_));
 OAI21_X1 _28902_ (.A(_02334_),
    .B1(_02336_),
    .B2(_02361_),
    .ZN(_03705_));
 OAI21_X1 _28903_ (.A(_02334_),
    .B1(_03062_),
    .B2(_02275_),
    .ZN(_03706_));
 AND4_X1 _28904_ (.A1(_03702_),
    .A2(_03704_),
    .A3(_03705_),
    .A4(_03706_),
    .ZN(_03707_));
 NAND4_X1 _28905_ (.A1(_03681_),
    .A2(_03693_),
    .A3(_03701_),
    .A4(_03707_),
    .ZN(_03708_));
 OAI211_X1 _28906_ (.A(_02369_),
    .B(_02162_),
    .C1(_02271_),
    .C2(_02301_),
    .ZN(_03709_));
 OAI21_X1 _28907_ (.A(_02369_),
    .B1(_02216_),
    .B2(_02309_),
    .ZN(_03710_));
 NAND3_X1 _28908_ (.A1(_03101_),
    .A2(_03709_),
    .A3(_03710_),
    .ZN(_03711_));
 OAI211_X1 _28909_ (.A(_02284_),
    .B(_02171_),
    .C1(_02288_),
    .C2(_02221_),
    .ZN(_03712_));
 OAI21_X1 _28910_ (.A(_03712_),
    .B1(_02373_),
    .B2(_03093_),
    .ZN(_03713_));
 AOI21_X1 _28911_ (.A(_03093_),
    .B1(_03462_),
    .B2(_02250_),
    .ZN(_03714_));
 AND2_X1 _28912_ (.A1(_02173_),
    .A2(_02317_),
    .ZN(_03715_));
 AND2_X1 _28913_ (.A1(_02173_),
    .A2(_02336_),
    .ZN(_03716_));
 OR2_X1 _28914_ (.A1(_03715_),
    .A2(_03716_),
    .ZN(_03717_));
 NOR4_X1 _28915_ (.A1(_03711_),
    .A2(_03713_),
    .A3(_03714_),
    .A4(_03717_),
    .ZN(_03718_));
 NAND2_X1 _28916_ (.A1(_02215_),
    .A2(_02159_),
    .ZN(_03719_));
 AND2_X1 _28917_ (.A1(_02209_),
    .A2(_02246_),
    .ZN(_03720_));
 NOR3_X1 _28918_ (.A1(_03106_),
    .A2(_03720_),
    .A3(_02322_),
    .ZN(_03721_));
 NAND2_X1 _28919_ (.A1(_02191_),
    .A2(_02317_),
    .ZN(_03722_));
 NAND4_X1 _28920_ (.A1(_02168_),
    .A2(_02157_),
    .A3(_02163_),
    .A4(_02178_),
    .ZN(_03723_));
 NAND4_X1 _28921_ (.A1(_02327_),
    .A2(_02168_),
    .A3(_02178_),
    .A4(_02259_),
    .ZN(_03724_));
 AND4_X1 _28922_ (.A1(_03722_),
    .A2(_03497_),
    .A3(_03723_),
    .A4(_03724_),
    .ZN(_03725_));
 OAI21_X1 _28923_ (.A(_02215_),
    .B1(_02200_),
    .B2(_02333_),
    .ZN(_03726_));
 AND4_X1 _28924_ (.A1(_03719_),
    .A2(_03721_),
    .A3(_03725_),
    .A4(_03726_),
    .ZN(_03728_));
 NAND2_X1 _28925_ (.A1(_02194_),
    .A2(_02351_),
    .ZN(_03729_));
 OAI21_X1 _28926_ (.A(_02325_),
    .B1(_02194_),
    .B2(_02204_),
    .ZN(_03730_));
 NAND2_X1 _28927_ (.A1(_02325_),
    .A2(_02356_),
    .ZN(_03731_));
 NAND2_X1 _28928_ (.A1(_02325_),
    .A2(_02268_),
    .ZN(_03732_));
 NAND2_X1 _28929_ (.A1(_02325_),
    .A2(_02278_),
    .ZN(_03733_));
 AND4_X1 _28930_ (.A1(_03730_),
    .A2(_03731_),
    .A3(_03732_),
    .A4(_03733_),
    .ZN(_03734_));
 OAI21_X1 _28931_ (.A(_02351_),
    .B1(_02328_),
    .B2(_02337_),
    .ZN(_03735_));
 OAI211_X1 _28932_ (.A(_02351_),
    .B(_02275_),
    .C1(_02188_),
    .C2(_02145_),
    .ZN(_03736_));
 AND4_X1 _28933_ (.A1(_03729_),
    .A2(_03734_),
    .A3(_03735_),
    .A4(_03736_),
    .ZN(_03737_));
 NAND2_X1 _28934_ (.A1(_02356_),
    .A2(_02358_),
    .ZN(_03739_));
 OAI21_X1 _28935_ (.A(_02180_),
    .B1(_02345_),
    .B2(_02311_),
    .ZN(_03740_));
 OAI21_X1 _28936_ (.A(_02292_),
    .B1(_03056_),
    .B2(_02336_),
    .ZN(_03741_));
 NAND2_X1 _28937_ (.A1(_02292_),
    .A2(_02199_),
    .ZN(_03742_));
 AND4_X1 _28938_ (.A1(_03739_),
    .A2(_03740_),
    .A3(_03741_),
    .A4(_03742_),
    .ZN(_03743_));
 NAND4_X1 _28939_ (.A1(_03718_),
    .A2(_03728_),
    .A3(_03737_),
    .A4(_03743_),
    .ZN(_03744_));
 NOR2_X1 _28940_ (.A1(_03708_),
    .A2(_03744_),
    .ZN(_03745_));
 INV_X1 _28941_ (.A(_03745_),
    .ZN(_03746_));
 XNOR2_X1 _28942_ (.A(_03670_),
    .B(_03746_),
    .ZN(_03747_));
 NAND3_X1 _28943_ (.A1(_03397_),
    .A2(_02061_),
    .A3(_01894_),
    .ZN(_03748_));
 OAI211_X1 _28944_ (.A(_03397_),
    .B(_01905_),
    .C1(_01954_),
    .C2(_03405_),
    .ZN(_03750_));
 OAI211_X1 _28945_ (.A(_03397_),
    .B(_01852_),
    .C1(_01856_),
    .C2(_01922_),
    .ZN(_03751_));
 OAI21_X1 _28946_ (.A(_03397_),
    .B1(_01945_),
    .B2(_01953_),
    .ZN(_03752_));
 AND4_X1 _28947_ (.A1(_03748_),
    .A2(_03750_),
    .A3(_03751_),
    .A4(_03752_),
    .ZN(_03753_));
 NAND4_X1 _28948_ (.A1(_01980_),
    .A2(_01846_),
    .A3(_01887_),
    .A4(_02103_),
    .ZN(_03754_));
 NAND4_X1 _28949_ (.A1(_01851_),
    .A2(_01980_),
    .A3(_01922_),
    .A4(_01887_),
    .ZN(_03755_));
 OAI211_X1 _28950_ (.A(_03754_),
    .B(_03755_),
    .C1(_02068_),
    .C2(_03386_),
    .ZN(_03756_));
 INV_X1 _28951_ (.A(_02042_),
    .ZN(_03757_));
 AOI21_X1 _28952_ (.A(_03386_),
    .B1(_02101_),
    .B2(_03757_),
    .ZN(_03758_));
 AND3_X1 _28953_ (.A1(_01882_),
    .A2(_01983_),
    .A3(_02072_),
    .ZN(_03759_));
 NOR3_X1 _28954_ (.A1(_03756_),
    .A2(_03758_),
    .A3(_03759_),
    .ZN(_03761_));
 AND2_X1 _28955_ (.A1(_02122_),
    .A2(_01901_),
    .ZN(_03762_));
 AND2_X1 _28956_ (.A1(_01973_),
    .A2(_01870_),
    .ZN(_03763_));
 NOR4_X1 _28957_ (.A1(_03762_),
    .A2(_03381_),
    .A3(_03763_),
    .A4(_02964_),
    .ZN(_03764_));
 OAI21_X1 _28958_ (.A(_01898_),
    .B1(_02971_),
    .B2(_02035_),
    .ZN(_03765_));
 NAND4_X1 _28959_ (.A1(_01851_),
    .A2(_01980_),
    .A3(_01922_),
    .A4(_01875_),
    .ZN(_03766_));
 AND3_X1 _28960_ (.A1(_03765_),
    .A2(_03378_),
    .A3(_03766_),
    .ZN(_03767_));
 AND2_X1 _28961_ (.A1(_02076_),
    .A2(_01961_),
    .ZN(_03768_));
 AND3_X1 _28962_ (.A1(_01884_),
    .A2(_02094_),
    .A3(_01896_),
    .ZN(_03769_));
 NOR4_X1 _28963_ (.A1(_03768_),
    .A2(_02981_),
    .A3(_03375_),
    .A4(_03769_),
    .ZN(_03770_));
 AND4_X1 _28964_ (.A1(_03761_),
    .A2(_03764_),
    .A3(_03767_),
    .A4(_03770_),
    .ZN(_03772_));
 OAI211_X1 _28965_ (.A(_03395_),
    .B(_02103_),
    .C1(_01894_),
    .C2(_01907_),
    .ZN(_03773_));
 OAI211_X1 _28966_ (.A(_03395_),
    .B(_01852_),
    .C1(_02088_),
    .C2(_01920_),
    .ZN(_03774_));
 OAI211_X1 _28967_ (.A(_03395_),
    .B(_01905_),
    .C1(_02088_),
    .C2(_03405_),
    .ZN(_03775_));
 OAI21_X1 _28968_ (.A(_03395_),
    .B1(_01979_),
    .B2(_03401_),
    .ZN(_03776_));
 AND4_X1 _28969_ (.A1(_03773_),
    .A2(_03774_),
    .A3(_03775_),
    .A4(_03776_),
    .ZN(_03777_));
 OAI21_X1 _28970_ (.A(_02059_),
    .B1(_01873_),
    .B2(_03442_),
    .ZN(_03778_));
 INV_X1 _28971_ (.A(_02023_),
    .ZN(_03779_));
 OAI21_X1 _28972_ (.A(_02059_),
    .B1(_03401_),
    .B2(_01903_),
    .ZN(_03780_));
 AND3_X1 _28973_ (.A1(_02052_),
    .A2(_03779_),
    .A3(_03780_),
    .ZN(_03781_));
 OAI21_X1 _28974_ (.A(_02031_),
    .B1(_02122_),
    .B2(_02108_),
    .ZN(_03783_));
 OAI21_X1 _28975_ (.A(_02031_),
    .B1(_01915_),
    .B2(_03401_),
    .ZN(_03784_));
 AND4_X1 _28976_ (.A1(_03778_),
    .A2(_03781_),
    .A3(_03783_),
    .A4(_03784_),
    .ZN(_03785_));
 AND4_X1 _28977_ (.A1(_03753_),
    .A2(_03772_),
    .A3(_03777_),
    .A4(_03785_),
    .ZN(_03786_));
 OAI21_X1 _28978_ (.A(_01843_),
    .B1(_01968_),
    .B2(_01915_),
    .ZN(_03787_));
 OAI21_X1 _28979_ (.A(_01843_),
    .B1(_02042_),
    .B2(_01963_),
    .ZN(_03788_));
 NAND3_X1 _28980_ (.A1(_02032_),
    .A2(_01885_),
    .A3(_01841_),
    .ZN(_03789_));
 AND4_X1 _28981_ (.A1(_03010_),
    .A2(_03787_),
    .A3(_03788_),
    .A4(_03789_),
    .ZN(_03790_));
 AND2_X1 _28982_ (.A1(_01867_),
    .A2(_01906_),
    .ZN(_03791_));
 OAI21_X1 _28983_ (.A(_01890_),
    .B1(_02042_),
    .B2(_03791_),
    .ZN(_03792_));
 NAND4_X1 _28984_ (.A1(_01935_),
    .A2(_03002_),
    .A3(_02009_),
    .A4(_01887_),
    .ZN(_03793_));
 AND4_X1 _28985_ (.A1(_01891_),
    .A2(_03790_),
    .A3(_03792_),
    .A4(_03793_),
    .ZN(_03794_));
 AOI21_X1 _28986_ (.A(_03431_),
    .B1(_01988_),
    .B2(_03426_),
    .ZN(_03795_));
 AOI21_X1 _28987_ (.A(_03795_),
    .B1(_01847_),
    .B2(_01992_),
    .ZN(_03796_));
 AND2_X1 _28988_ (.A1(_01979_),
    .A2(_01958_),
    .ZN(_03797_));
 AOI211_X1 _28989_ (.A(_03797_),
    .B(_02119_),
    .C1(_01915_),
    .C2(_01992_),
    .ZN(_03798_));
 OAI21_X1 _28990_ (.A(_01952_),
    .B1(_01945_),
    .B2(_01953_),
    .ZN(_03799_));
 NAND2_X1 _28991_ (.A1(_01952_),
    .A2(_01949_),
    .ZN(_03800_));
 AND2_X1 _28992_ (.A1(_03799_),
    .A2(_03800_),
    .ZN(_03801_));
 OAI21_X1 _28993_ (.A(_01952_),
    .B1(_01996_),
    .B2(_01979_),
    .ZN(_03802_));
 AND4_X1 _28994_ (.A1(_03796_),
    .A2(_03798_),
    .A3(_03801_),
    .A4(_03802_),
    .ZN(_03804_));
 AOI211_X1 _28995_ (.A(_01927_),
    .B(_01879_),
    .C1(_02088_),
    .C2(_03405_),
    .ZN(_03805_));
 OAI21_X1 _28996_ (.A(_01855_),
    .B1(_01963_),
    .B2(_01902_),
    .ZN(_03806_));
 OAI211_X1 _28997_ (.A(_03002_),
    .B(_03003_),
    .C1(_01884_),
    .C2(_01858_),
    .ZN(_03807_));
 NAND2_X1 _28998_ (.A1(_02014_),
    .A2(_02035_),
    .ZN(_03808_));
 NAND4_X1 _28999_ (.A1(_03806_),
    .A2(_03807_),
    .A3(_03007_),
    .A4(_03808_),
    .ZN(_03809_));
 AND2_X1 _29000_ (.A1(_02986_),
    .A2(_02047_),
    .ZN(_03810_));
 INV_X1 _29001_ (.A(_01939_),
    .ZN(_03811_));
 AOI21_X1 _29002_ (.A(_01879_),
    .B1(_01969_),
    .B2(_03811_),
    .ZN(_03812_));
 NOR4_X1 _29003_ (.A1(_03805_),
    .A2(_03809_),
    .A3(_03810_),
    .A4(_03812_),
    .ZN(_03813_));
 NAND2_X1 _29004_ (.A1(_01979_),
    .A2(_02132_),
    .ZN(_03815_));
 OAI21_X1 _29005_ (.A(_01934_),
    .B1(_02108_),
    .B2(_01884_),
    .ZN(_03816_));
 NAND3_X1 _29006_ (.A1(_01895_),
    .A2(_02072_),
    .A3(_02132_),
    .ZN(_03817_));
 NAND2_X1 _29007_ (.A1(_01934_),
    .A2(_02042_),
    .ZN(_03818_));
 AND4_X1 _29008_ (.A1(_03815_),
    .A2(_03816_),
    .A3(_03817_),
    .A4(_03818_),
    .ZN(_03819_));
 AND4_X1 _29009_ (.A1(_03794_),
    .A2(_03804_),
    .A3(_03813_),
    .A4(_03819_),
    .ZN(_03820_));
 NAND2_X2 _29010_ (.A1(_03786_),
    .A2(_03820_),
    .ZN(_03821_));
 INV_X1 _29011_ (.A(_02533_),
    .ZN(_03822_));
 INV_X1 _29012_ (.A(_02610_),
    .ZN(_03823_));
 OAI21_X1 _29013_ (.A(_03318_),
    .B1(_03822_),
    .B2(_03823_),
    .ZN(_03824_));
 AND2_X1 _29014_ (.A1(_02921_),
    .A2(_02534_),
    .ZN(_03826_));
 AOI211_X1 _29015_ (.A(_03824_),
    .B(_03826_),
    .C1(_02454_),
    .C2(_02534_),
    .ZN(_03827_));
 OAI21_X1 _29016_ (.A(_02561_),
    .B1(_03324_),
    .B2(_02468_),
    .ZN(_03828_));
 NAND4_X1 _29017_ (.A1(_03322_),
    .A2(_02553_),
    .A3(_02452_),
    .A4(_02558_),
    .ZN(_03829_));
 AND3_X1 _29018_ (.A1(_03828_),
    .A2(_03314_),
    .A3(_03829_),
    .ZN(_03830_));
 OAI211_X1 _29019_ (.A(_02549_),
    .B(_02435_),
    .C1(_02452_),
    .C2(_02423_),
    .ZN(_03831_));
 INV_X1 _29020_ (.A(_02523_),
    .ZN(_03832_));
 OAI211_X1 _29021_ (.A(_03831_),
    .B(_02940_),
    .C1(_03832_),
    .C2(_02938_),
    .ZN(_03833_));
 AND4_X1 _29022_ (.A1(_02429_),
    .A2(_02553_),
    .A3(_02470_),
    .A4(_02554_),
    .ZN(_03834_));
 AOI21_X1 _29023_ (.A(_02938_),
    .B1(_02544_),
    .B2(_03367_),
    .ZN(_03835_));
 NOR3_X1 _29024_ (.A1(_03833_),
    .A2(_03834_),
    .A3(_03835_),
    .ZN(_03837_));
 AND2_X1 _29025_ (.A1(_02537_),
    .A2(_02458_),
    .ZN(_03838_));
 AND2_X1 _29026_ (.A1(_02537_),
    .A2(_02924_),
    .ZN(_03839_));
 NOR2_X1 _29027_ (.A1(_03838_),
    .A2(_03839_),
    .ZN(_03840_));
 AND4_X1 _29028_ (.A1(_02539_),
    .A2(_03840_),
    .A3(_02955_),
    .A4(_03321_),
    .ZN(_03841_));
 NAND4_X1 _29029_ (.A1(_03827_),
    .A2(_03830_),
    .A3(_03837_),
    .A4(_03841_),
    .ZN(_03842_));
 OAI211_X1 _29030_ (.A(_02441_),
    .B(_02470_),
    .C1(_02472_),
    .C2(_02397_),
    .ZN(_03843_));
 OAI211_X1 _29031_ (.A(_02441_),
    .B(_02394_),
    .C1(_02880_),
    .C2(_02557_),
    .ZN(_03844_));
 OAI211_X1 _29032_ (.A(_02441_),
    .B(_02435_),
    .C1(_02880_),
    .C2(_02429_),
    .ZN(_03845_));
 OAI21_X1 _29033_ (.A(_02441_),
    .B1(_02527_),
    .B2(_02522_),
    .ZN(_03846_));
 AND4_X1 _29034_ (.A1(_03843_),
    .A2(_03844_),
    .A3(_03845_),
    .A4(_03846_),
    .ZN(_03848_));
 NAND2_X1 _29035_ (.A1(_02420_),
    .A2(_02461_),
    .ZN(_03849_));
 NAND2_X1 _29036_ (.A1(_02468_),
    .A2(_02461_),
    .ZN(_03850_));
 AND3_X1 _29037_ (.A1(_03849_),
    .A2(_03850_),
    .A3(_02473_),
    .ZN(_03851_));
 OAI21_X1 _29038_ (.A(_02462_),
    .B1(_02446_),
    .B2(_02495_),
    .ZN(_03852_));
 OAI211_X1 _29039_ (.A(_02462_),
    .B(_03322_),
    .C1(_02452_),
    .C2(_02423_),
    .ZN(_03853_));
 NAND4_X1 _29040_ (.A1(_03848_),
    .A2(_03851_),
    .A3(_03852_),
    .A4(_03853_),
    .ZN(_03854_));
 OAI21_X1 _29041_ (.A(_02432_),
    .B1(_02541_),
    .B2(_02523_),
    .ZN(_03855_));
 OAI211_X1 _29042_ (.A(_02432_),
    .B(_02435_),
    .C1(_02880_),
    .C2(_02430_),
    .ZN(_03856_));
 OAI21_X1 _29043_ (.A(_02432_),
    .B1(_02578_),
    .B2(_02571_),
    .ZN(_03857_));
 NAND4_X1 _29044_ (.A1(_03322_),
    .A2(_02438_),
    .A3(_02452_),
    .A4(_02558_),
    .ZN(_03858_));
 NAND4_X1 _29045_ (.A1(_03855_),
    .A2(_03856_),
    .A3(_03857_),
    .A4(_03858_),
    .ZN(_03859_));
 AND3_X1 _29046_ (.A1(_02602_),
    .A2(_03295_),
    .A3(_02438_),
    .ZN(_03860_));
 AND3_X1 _29047_ (.A1(_02547_),
    .A2(_02391_),
    .A3(_02927_),
    .ZN(_03861_));
 AND2_X1 _29048_ (.A1(_02391_),
    .A2(_02424_),
    .ZN(_03862_));
 OR4_X1 _29049_ (.A1(_03860_),
    .A2(_03861_),
    .A3(_03291_),
    .A4(_03862_),
    .ZN(_03863_));
 NOR4_X1 _29050_ (.A1(_03842_),
    .A2(_03854_),
    .A3(_03859_),
    .A4(_03863_),
    .ZN(_03864_));
 NAND2_X1 _29051_ (.A1(_02504_),
    .A2(_02450_),
    .ZN(_03865_));
 OAI21_X1 _29052_ (.A(_02503_),
    .B1(_02446_),
    .B2(_02495_),
    .ZN(_03866_));
 NAND3_X1 _29053_ (.A1(_02527_),
    .A2(_03295_),
    .A3(_02524_),
    .ZN(_03867_));
 AND4_X1 _29054_ (.A1(_02505_),
    .A2(_03865_),
    .A3(_03866_),
    .A4(_03867_),
    .ZN(_03869_));
 NAND4_X1 _29055_ (.A1(_02470_),
    .A2(_02558_),
    .A3(_02524_),
    .A4(_02430_),
    .ZN(_03870_));
 OAI211_X1 _29056_ (.A(_02498_),
    .B(_03322_),
    .C1(_02472_),
    .C2(_02397_),
    .ZN(_03871_));
 AND2_X1 _29057_ (.A1(_02527_),
    .A2(_02493_),
    .ZN(_03872_));
 AND3_X1 _29058_ (.A1(_02493_),
    .A2(_02472_),
    .A3(_02454_),
    .ZN(_03873_));
 AOI211_X1 _29059_ (.A(_03872_),
    .B(_03873_),
    .C1(_02595_),
    .C2(_02498_),
    .ZN(_03874_));
 NAND4_X1 _29060_ (.A1(_03869_),
    .A2(_03870_),
    .A3(_03871_),
    .A4(_03874_),
    .ZN(_03875_));
 OAI211_X1 _29061_ (.A(_02586_),
    .B(_02583_),
    .C1(_02610_),
    .C2(_02443_),
    .ZN(_03876_));
 NAND2_X1 _29062_ (.A1(_02574_),
    .A2(_02454_),
    .ZN(_03877_));
 NAND2_X1 _29063_ (.A1(_02574_),
    .A2(_02467_),
    .ZN(_03878_));
 NAND4_X1 _29064_ (.A1(_03876_),
    .A2(_02929_),
    .A3(_03877_),
    .A4(_03878_),
    .ZN(_03880_));
 AOI21_X1 _29065_ (.A(_02569_),
    .B1(_02447_),
    .B2(_03297_),
    .ZN(_03881_));
 AND2_X1 _29066_ (.A1(_02407_),
    .A2(_02395_),
    .ZN(_03882_));
 INV_X1 _29067_ (.A(_03882_),
    .ZN(_03883_));
 AOI21_X1 _29068_ (.A(_02569_),
    .B1(_02421_),
    .B2(_03883_),
    .ZN(_03884_));
 OR4_X1 _29069_ (.A1(_02913_),
    .A2(_03880_),
    .A3(_03881_),
    .A4(_03884_),
    .ZN(_03885_));
 OAI21_X1 _29070_ (.A(_02593_),
    .B1(_02509_),
    .B2(_02578_),
    .ZN(_03886_));
 OAI21_X1 _29071_ (.A(_02600_),
    .B1(_02563_),
    .B2(_02564_),
    .ZN(_03887_));
 AND2_X1 _29072_ (.A1(_02434_),
    .A2(_02557_),
    .ZN(_03888_));
 OAI21_X1 _29073_ (.A(_02593_),
    .B1(_02408_),
    .B2(_03888_),
    .ZN(_03889_));
 OAI21_X1 _29074_ (.A(_02599_),
    .B1(_02398_),
    .B2(_02486_),
    .ZN(_03891_));
 NAND4_X1 _29075_ (.A1(_03886_),
    .A2(_03887_),
    .A3(_03889_),
    .A4(_03891_),
    .ZN(_03892_));
 AND2_X1 _29076_ (.A1(_02527_),
    .A2(_02479_),
    .ZN(_03893_));
 INV_X1 _29077_ (.A(_02924_),
    .ZN(_03894_));
 NAND2_X1 _29078_ (.A1(_02544_),
    .A2(_03894_),
    .ZN(_03895_));
 AOI21_X1 _29079_ (.A(_03893_),
    .B1(_03895_),
    .B2(_02479_),
    .ZN(_03896_));
 NAND2_X1 _29080_ (.A1(_02515_),
    .A2(_02610_),
    .ZN(_03897_));
 NAND2_X1 _29081_ (.A1(_02602_),
    .A2(_02515_),
    .ZN(_03898_));
 NAND2_X1 _29082_ (.A1(_02514_),
    .A2(_02408_),
    .ZN(_03899_));
 NAND4_X1 _29083_ (.A1(_03896_),
    .A2(_03897_),
    .A3(_03898_),
    .A4(_03899_),
    .ZN(_03900_));
 NOR4_X1 _29084_ (.A1(_03875_),
    .A2(_03885_),
    .A3(_03892_),
    .A4(_03900_),
    .ZN(_03901_));
 NAND2_X2 _29085_ (.A1(_03864_),
    .A2(_03901_),
    .ZN(_03902_));
 XOR2_X1 _29086_ (.A(_03821_),
    .B(_03902_),
    .Z(_03903_));
 OAI21_X1 _29087_ (.A(_02759_),
    .B1(_02727_),
    .B2(_02728_),
    .ZN(_03904_));
 NAND4_X1 _29088_ (.A1(_02759_),
    .A2(_02775_),
    .A3(_02667_),
    .A4(_02832_),
    .ZN(_03905_));
 NAND4_X1 _29089_ (.A1(_03904_),
    .A2(_03905_),
    .A3(_03177_),
    .A4(_03567_),
    .ZN(_03906_));
 AND2_X1 _29090_ (.A1(_02764_),
    .A2(_02728_),
    .ZN(_03907_));
 NOR2_X1 _29091_ (.A1(_03907_),
    .A2(_02766_),
    .ZN(_03908_));
 OAI21_X1 _29092_ (.A(_03908_),
    .B1(_02772_),
    .B2(_02719_),
    .ZN(_03909_));
 AOI211_X1 _29093_ (.A(_03906_),
    .B(_03909_),
    .C1(_03172_),
    .C2(_02737_),
    .ZN(_03910_));
 NAND2_X1 _29094_ (.A1(_02832_),
    .A2(_02666_),
    .ZN(_03912_));
 INV_X1 _29095_ (.A(_03912_),
    .ZN(_03913_));
 NAND2_X1 _29096_ (.A1(_03913_),
    .A2(_02811_),
    .ZN(_03914_));
 AND2_X1 _29097_ (.A1(_02805_),
    .A2(_02796_),
    .ZN(_03915_));
 AND2_X1 _29098_ (.A1(_02805_),
    .A2(_02675_),
    .ZN(_03916_));
 AND2_X1 _29099_ (.A1(_02805_),
    .A2(_03156_),
    .ZN(_03917_));
 NOR4_X1 _29100_ (.A1(_03915_),
    .A2(_03916_),
    .A3(_03917_),
    .A4(_03608_),
    .ZN(_03918_));
 NAND2_X1 _29101_ (.A1(_02812_),
    .A2(_03246_),
    .ZN(_03919_));
 OAI211_X1 _29102_ (.A(_02812_),
    .B(_16778_),
    .C1(_02657_),
    .C2(_02650_),
    .ZN(_03920_));
 AND4_X1 _29103_ (.A1(_03914_),
    .A2(_03918_),
    .A3(_03919_),
    .A4(_03920_),
    .ZN(_03921_));
 OAI211_X1 _29104_ (.A(_03204_),
    .B(_03549_),
    .C1(_02747_),
    .C2(_02642_),
    .ZN(_03923_));
 NAND2_X1 _29105_ (.A1(_02789_),
    .A2(_03923_),
    .ZN(_03924_));
 OAI211_X1 _29106_ (.A(_02799_),
    .B(_03549_),
    .C1(_02638_),
    .C2(_03528_),
    .ZN(_03925_));
 OAI21_X1 _29107_ (.A(_02799_),
    .B1(_02724_),
    .B2(_03156_),
    .ZN(_03926_));
 OAI21_X1 _29108_ (.A(_02799_),
    .B1(_02765_),
    .B2(_02671_),
    .ZN(_03927_));
 NAND2_X1 _29109_ (.A1(_02799_),
    .A2(_02737_),
    .ZN(_03928_));
 NAND4_X1 _29110_ (.A1(_03925_),
    .A2(_03926_),
    .A3(_03927_),
    .A4(_03928_),
    .ZN(_03929_));
 AOI21_X1 _29111_ (.A(_03190_),
    .B1(_02773_),
    .B2(_02816_),
    .ZN(_03930_));
 NOR4_X1 _29112_ (.A1(_03924_),
    .A2(_03929_),
    .A3(_02792_),
    .A4(_03930_),
    .ZN(_03931_));
 OAI211_X1 _29113_ (.A(_02828_),
    .B(_03246_),
    .C1(_02747_),
    .C2(_02642_),
    .ZN(_03932_));
 NAND2_X1 _29114_ (.A1(_03558_),
    .A2(_02821_),
    .ZN(_03934_));
 OAI211_X1 _29115_ (.A(_03932_),
    .B(_03934_),
    .C1(_03193_),
    .C2(_03151_),
    .ZN(_03935_));
 NAND2_X1 _29116_ (.A1(_02831_),
    .A2(_02658_),
    .ZN(_03936_));
 OAI211_X1 _29117_ (.A(_03936_),
    .B(_03601_),
    .C1(_03229_),
    .C2(_03189_),
    .ZN(_03937_));
 AOI21_X1 _29118_ (.A(_03189_),
    .B1(_02808_),
    .B2(_03572_),
    .ZN(_03938_));
 NAND4_X1 _29119_ (.A1(_03211_),
    .A2(_03528_),
    .A3(_02702_),
    .A4(_03234_),
    .ZN(_03939_));
 OAI21_X1 _29120_ (.A(_03939_),
    .B1(_03189_),
    .B2(_03207_),
    .ZN(_03940_));
 NOR4_X1 _29121_ (.A1(_03935_),
    .A2(_03937_),
    .A3(_03938_),
    .A4(_03940_),
    .ZN(_03941_));
 AND4_X1 _29122_ (.A1(_03910_),
    .A2(_03921_),
    .A3(_03931_),
    .A4(_03941_),
    .ZN(_03942_));
 AND2_X1 _29123_ (.A1(_02664_),
    .A2(_02711_),
    .ZN(_03943_));
 INV_X1 _29124_ (.A(_03943_),
    .ZN(_03945_));
 NAND2_X1 _29125_ (.A1(_02665_),
    .A2(_02724_),
    .ZN(_03946_));
 OAI211_X1 _29126_ (.A(_03945_),
    .B(_03946_),
    .C1(_03581_),
    .C2(_02688_),
    .ZN(_03947_));
 NAND2_X1 _29127_ (.A1(_03148_),
    .A2(_03549_),
    .ZN(_03948_));
 AOI21_X1 _29128_ (.A(_03581_),
    .B1(_03151_),
    .B2(_03948_),
    .ZN(_03949_));
 INV_X1 _29129_ (.A(_02635_),
    .ZN(_03950_));
 AOI21_X1 _29130_ (.A(_03950_),
    .B1(_03571_),
    .B2(_03207_),
    .ZN(_03951_));
 BUF_X2 _29131_ (.A(_02815_),
    .Z(_03952_));
 NAND2_X1 _29132_ (.A1(_02635_),
    .A2(_03952_),
    .ZN(_03953_));
 NAND2_X1 _29133_ (.A1(_03210_),
    .A2(_03953_),
    .ZN(_03954_));
 NOR4_X1 _29134_ (.A1(_03947_),
    .A2(_03949_),
    .A3(_03951_),
    .A4(_03954_),
    .ZN(_03956_));
 OAI21_X1 _29135_ (.A(_02733_),
    .B1(_03160_),
    .B2(_02696_),
    .ZN(_03957_));
 AND4_X1 _29136_ (.A1(_02800_),
    .A2(_02662_),
    .A3(_02652_),
    .A4(_02678_),
    .ZN(_03958_));
 AND4_X1 _29137_ (.A1(_02662_),
    .A2(_02627_),
    .A3(_02702_),
    .A4(_02678_),
    .ZN(_03959_));
 AOI211_X1 _29138_ (.A(_03958_),
    .B(_03959_),
    .C1(_02813_),
    .C2(_02742_),
    .ZN(_03960_));
 OAI21_X1 _29139_ (.A(_02733_),
    .B1(_03182_),
    .B2(_02728_),
    .ZN(_03961_));
 NAND2_X1 _29140_ (.A1(_02742_),
    .A2(_02658_),
    .ZN(_03962_));
 AND4_X1 _29141_ (.A1(_02738_),
    .A2(_03962_),
    .A3(_03538_),
    .A4(_02740_),
    .ZN(_03963_));
 AND4_X1 _29142_ (.A1(_03957_),
    .A2(_03960_),
    .A3(_03961_),
    .A4(_03963_),
    .ZN(_03964_));
 OAI21_X1 _29143_ (.A(_02723_),
    .B1(_02711_),
    .B2(_02698_),
    .ZN(_03965_));
 OAI21_X1 _29144_ (.A(_02723_),
    .B1(_03558_),
    .B2(_02671_),
    .ZN(_03967_));
 OAI21_X1 _29145_ (.A(_02717_),
    .B1(_02711_),
    .B2(_03952_),
    .ZN(_03968_));
 OAI21_X1 _29146_ (.A(_02717_),
    .B1(_03558_),
    .B2(_02728_),
    .ZN(_03969_));
 AND4_X1 _29147_ (.A1(_03965_),
    .A2(_03967_),
    .A3(_03968_),
    .A4(_03969_),
    .ZN(_03970_));
 NAND2_X1 _29148_ (.A1(_03532_),
    .A2(_02832_),
    .ZN(_03971_));
 NAND3_X1 _29149_ (.A1(_03175_),
    .A2(_03528_),
    .A3(_03549_),
    .ZN(_03972_));
 NAND2_X1 _29150_ (.A1(_03971_),
    .A2(_03972_),
    .ZN(_03973_));
 OAI211_X1 _29151_ (.A(_03541_),
    .B(_03549_),
    .C1(_02747_),
    .C2(_02657_),
    .ZN(_03974_));
 OAI21_X1 _29152_ (.A(_03541_),
    .B1(_02782_),
    .B2(_03952_),
    .ZN(_03975_));
 NAND3_X1 _29153_ (.A1(_03974_),
    .A2(_03975_),
    .A3(_02706_),
    .ZN(_03976_));
 AND2_X1 _29154_ (.A1(_02737_),
    .A2(_03175_),
    .ZN(_03978_));
 NOR2_X1 _29155_ (.A1(_02691_),
    .A2(_03201_),
    .ZN(_03979_));
 NOR4_X1 _29156_ (.A1(_03973_),
    .A2(_03976_),
    .A3(_03978_),
    .A4(_03979_),
    .ZN(_03980_));
 AND4_X1 _29157_ (.A1(_03956_),
    .A2(_03964_),
    .A3(_03970_),
    .A4(_03980_),
    .ZN(_03981_));
 NAND2_X2 _29158_ (.A1(_03942_),
    .A2(_03981_),
    .ZN(_03982_));
 XOR2_X1 _29159_ (.A(_03982_),
    .B(_02837_),
    .Z(_03983_));
 XNOR2_X1 _29160_ (.A(_03903_),
    .B(_03983_),
    .ZN(_03984_));
 XNOR2_X1 _29161_ (.A(_03747_),
    .B(_03984_),
    .ZN(_03985_));
 XNOR2_X1 _29162_ (.A(_03985_),
    .B(_17156_),
    .ZN(_03986_));
 MUX2_X1 _29163_ (.A(_03669_),
    .B(_03986_),
    .S(_01825_),
    .Z(_00711_));
 XOR2_X1 _29164_ (.A(_17157_),
    .B(_17027_),
    .Z(_03987_));
 XOR2_X2 _29165_ (.A(_02139_),
    .B(_03821_),
    .Z(_03988_));
 OAI211_X1 _29166_ (.A(_02284_),
    .B(_02178_),
    .C1(_02223_),
    .C2(_02333_),
    .ZN(_03989_));
 OAI21_X1 _29167_ (.A(_02215_),
    .B1(_03118_),
    .B2(_02363_),
    .ZN(_03990_));
 OAI21_X1 _29168_ (.A(_02215_),
    .B1(_02200_),
    .B2(_02356_),
    .ZN(_03991_));
 AND4_X1 _29169_ (.A1(_03719_),
    .A2(_03990_),
    .A3(_02343_),
    .A4(_03991_),
    .ZN(_03992_));
 NAND2_X1 _29170_ (.A1(_02191_),
    .A2(_03061_),
    .ZN(_03993_));
 OAI211_X1 _29171_ (.A(_02284_),
    .B(_02178_),
    .C1(_02347_),
    .C2(_02353_),
    .ZN(_03994_));
 AND4_X1 _29172_ (.A1(_03989_),
    .A2(_03992_),
    .A3(_03993_),
    .A4(_03994_),
    .ZN(_03995_));
 AND2_X1 _29173_ (.A1(_02212_),
    .A2(_02370_),
    .ZN(_03996_));
 AND2_X1 _29174_ (.A1(_02173_),
    .A2(_02246_),
    .ZN(_03998_));
 AOI211_X1 _29175_ (.A(_03996_),
    .B(_03998_),
    .C1(_02368_),
    .C2(_02212_),
    .ZN(_03999_));
 AND3_X1 _29176_ (.A1(_02363_),
    .A2(_02284_),
    .A3(_02150_),
    .ZN(_04000_));
 AOI211_X1 _29177_ (.A(_04000_),
    .B(_02316_),
    .C1(_02369_),
    .C2(_02318_),
    .ZN(_04001_));
 OAI21_X1 _29178_ (.A(_02212_),
    .B1(_02288_),
    .B2(_02379_),
    .ZN(_04002_));
 AND4_X1 _29179_ (.A1(_03103_),
    .A2(_03999_),
    .A3(_04001_),
    .A4(_04002_),
    .ZN(_04003_));
 NAND2_X1 _29180_ (.A1(_02176_),
    .A2(_02380_),
    .ZN(_04004_));
 NAND3_X1 _29181_ (.A1(_02380_),
    .A2(_02352_),
    .A3(_02145_),
    .ZN(_04005_));
 NAND4_X1 _29182_ (.A1(_04004_),
    .A2(_03071_),
    .A3(_03502_),
    .A4(_04005_),
    .ZN(_04006_));
 NAND2_X1 _29183_ (.A1(_02325_),
    .A2(_02216_),
    .ZN(_04007_));
 NAND3_X1 _29184_ (.A1(_04007_),
    .A2(_03731_),
    .A3(_03079_),
    .ZN(_04008_));
 AND2_X1 _29185_ (.A1(_02326_),
    .A2(_02318_),
    .ZN(_04009_));
 AND2_X1 _29186_ (.A1(_02189_),
    .A2(_02326_),
    .ZN(_04010_));
 NOR4_X1 _29187_ (.A1(_04006_),
    .A2(_04008_),
    .A3(_04009_),
    .A4(_04010_),
    .ZN(_04011_));
 NAND3_X1 _29188_ (.A1(_02231_),
    .A2(_02239_),
    .A3(_02339_),
    .ZN(_04012_));
 AND2_X1 _29189_ (.A1(_02332_),
    .A2(_02180_),
    .ZN(_04013_));
 AND3_X1 _29190_ (.A1(_02358_),
    .A2(_02198_),
    .A3(_02225_),
    .ZN(_04014_));
 AOI211_X1 _29191_ (.A(_04013_),
    .B(_04014_),
    .C1(_02358_),
    .C2(_02189_),
    .ZN(_04015_));
 OAI211_X1 _29192_ (.A(_02339_),
    .B(_02259_),
    .C1(_02162_),
    .C2(_02353_),
    .ZN(_04016_));
 OAI21_X1 _29193_ (.A(_02339_),
    .B1(_02223_),
    .B2(_02333_),
    .ZN(_04017_));
 AND4_X1 _29194_ (.A1(_04012_),
    .A2(_04015_),
    .A3(_04016_),
    .A4(_04017_),
    .ZN(_04019_));
 NAND4_X1 _29195_ (.A1(_03995_),
    .A2(_04003_),
    .A3(_04011_),
    .A4(_04019_),
    .ZN(_04020_));
 INV_X1 _29196_ (.A(_02229_),
    .ZN(_04021_));
 AND2_X1 _29197_ (.A1(_02220_),
    .A2(_02247_),
    .ZN(_04022_));
 AOI211_X1 _29198_ (.A(_03674_),
    .B(_04022_),
    .C1(_03056_),
    .C2(_02220_),
    .ZN(_04023_));
 OAI21_X1 _29199_ (.A(_03052_),
    .B1(_02246_),
    .B2(_02248_),
    .ZN(_04024_));
 OAI21_X1 _29200_ (.A(_03052_),
    .B1(_03062_),
    .B2(_02200_),
    .ZN(_04025_));
 AND4_X1 _29201_ (.A1(_04021_),
    .A2(_04023_),
    .A3(_04024_),
    .A4(_04025_),
    .ZN(_04026_));
 INV_X1 _29202_ (.A(_02312_),
    .ZN(_04027_));
 OAI21_X1 _29203_ (.A(_02235_),
    .B1(_02176_),
    .B2(_02336_),
    .ZN(_04028_));
 OAI211_X1 _29204_ (.A(_02308_),
    .B(_16770_),
    .C1(_16769_),
    .C2(_02198_),
    .ZN(_04029_));
 OAI21_X1 _29205_ (.A(_02235_),
    .B1(_02252_),
    .B2(_02276_),
    .ZN(_04030_));
 AND4_X1 _29206_ (.A1(_04027_),
    .A2(_04028_),
    .A3(_04029_),
    .A4(_04030_),
    .ZN(_04031_));
 AND2_X1 _29207_ (.A1(_02244_),
    .A2(_02320_),
    .ZN(_04032_));
 INV_X1 _29208_ (.A(_04032_),
    .ZN(_04033_));
 OAI21_X1 _29209_ (.A(_02245_),
    .B1(_02248_),
    .B2(_02370_),
    .ZN(_04034_));
 OAI211_X1 _29210_ (.A(_02245_),
    .B(_02352_),
    .C1(_03075_),
    .C2(_02285_),
    .ZN(_04035_));
 NAND4_X1 _29211_ (.A1(_04033_),
    .A2(_03698_),
    .A3(_04034_),
    .A4(_04035_),
    .ZN(_04036_));
 AND2_X1 _29212_ (.A1(_02264_),
    .A2(_02370_),
    .ZN(_04037_));
 AND2_X1 _29213_ (.A1(_03081_),
    .A2(_02265_),
    .ZN(_04038_));
 NOR4_X1 _29214_ (.A1(_04036_),
    .A2(_04037_),
    .A3(_04038_),
    .A4(_03474_),
    .ZN(_04040_));
 AOI22_X1 _29215_ (.A1(_03064_),
    .A2(_02239_),
    .B1(_02379_),
    .B2(_02334_),
    .ZN(_04041_));
 OAI21_X1 _29216_ (.A(_02334_),
    .B1(_02363_),
    .B2(_02318_),
    .ZN(_04042_));
 OAI21_X1 _29217_ (.A(_02152_),
    .B1(_02146_),
    .B2(_02379_),
    .ZN(_04043_));
 AND4_X1 _29218_ (.A1(_03046_),
    .A2(_04041_),
    .A3(_04042_),
    .A4(_04043_),
    .ZN(_04044_));
 NAND4_X1 _29219_ (.A1(_04026_),
    .A2(_04031_),
    .A3(_04040_),
    .A4(_04044_),
    .ZN(_04045_));
 NOR2_X2 _29220_ (.A1(_04020_),
    .A2(_04045_),
    .ZN(_04046_));
 XNOR2_X1 _29221_ (.A(_03988_),
    .B(_04046_),
    .ZN(_04047_));
 NAND2_X1 _29222_ (.A1(_02686_),
    .A2(_03204_),
    .ZN(_04048_));
 NAND2_X1 _29223_ (.A1(_02780_),
    .A2(_02643_),
    .ZN(_04049_));
 NAND2_X1 _29224_ (.A1(_02798_),
    .A2(_04049_),
    .ZN(_04050_));
 AND2_X1 _29225_ (.A1(_02780_),
    .A2(_02696_),
    .ZN(_04051_));
 AOI221_X1 _29226_ (.A(_04050_),
    .B1(_02626_),
    .B2(_04051_),
    .C1(_02799_),
    .C2(_02689_),
    .ZN(_04052_));
 OAI21_X1 _29227_ (.A(_03204_),
    .B1(_03952_),
    .B2(_02696_),
    .ZN(_04053_));
 NOR4_X1 _29228_ (.A1(_03555_),
    .A2(_02786_),
    .A3(_02790_),
    .A4(_03215_),
    .ZN(_04054_));
 AND4_X1 _29229_ (.A1(_04048_),
    .A2(_04052_),
    .A3(_04053_),
    .A4(_04054_),
    .ZN(_04055_));
 OAI21_X1 _29230_ (.A(_02754_),
    .B1(_02689_),
    .B2(_03230_),
    .ZN(_04056_));
 INV_X1 _29231_ (.A(_03221_),
    .ZN(_04057_));
 NAND3_X1 _29232_ (.A1(_02754_),
    .A2(_02800_),
    .A3(_03528_),
    .ZN(_04058_));
 AND4_X1 _29233_ (.A1(_02756_),
    .A2(_04056_),
    .A3(_04057_),
    .A4(_04058_),
    .ZN(_04059_));
 OAI21_X1 _29234_ (.A(_02769_),
    .B1(_02711_),
    .B2(_02686_),
    .ZN(_04060_));
 OAI211_X1 _29235_ (.A(_02769_),
    .B(_02667_),
    .C1(_02638_),
    .C2(_03528_),
    .ZN(_04061_));
 NAND2_X1 _29236_ (.A1(_02782_),
    .A2(_02769_),
    .ZN(_04062_));
 AND3_X1 _29237_ (.A1(_04060_),
    .A2(_04061_),
    .A3(_04062_),
    .ZN(_04063_));
 OAI211_X1 _29238_ (.A(_03172_),
    .B(_03549_),
    .C1(_02747_),
    .C2(_02657_),
    .ZN(_04064_));
 OAI21_X1 _29239_ (.A(_03172_),
    .B1(_02765_),
    .B2(_02671_),
    .ZN(_04065_));
 AND4_X1 _29240_ (.A1(_04059_),
    .A2(_04063_),
    .A3(_04064_),
    .A4(_04065_),
    .ZN(_04066_));
 OAI21_X1 _29241_ (.A(_02812_),
    .B1(_03913_),
    .B2(_02686_),
    .ZN(_04067_));
 AOI21_X1 _29242_ (.A(_03607_),
    .B1(_02720_),
    .B2(_02805_),
    .ZN(_04068_));
 OAI21_X1 _29243_ (.A(_02812_),
    .B1(_03150_),
    .B2(_02727_),
    .ZN(_04069_));
 OAI21_X1 _29244_ (.A(_02805_),
    .B1(_03209_),
    .B2(_03156_),
    .ZN(_04070_));
 AND4_X1 _29245_ (.A1(_04067_),
    .A2(_04068_),
    .A3(_04069_),
    .A4(_04070_),
    .ZN(_04071_));
 AND2_X1 _29246_ (.A1(_02821_),
    .A2(_02686_),
    .ZN(_04072_));
 AND2_X1 _29247_ (.A1(_02821_),
    .A2(_02654_),
    .ZN(_04073_));
 NOR2_X1 _29248_ (.A1(_04072_),
    .A2(_04073_),
    .ZN(_04074_));
 OAI21_X1 _29249_ (.A(_02828_),
    .B1(_03558_),
    .B2(_02704_),
    .ZN(_04075_));
 OAI211_X1 _29250_ (.A(_04074_),
    .B(_04075_),
    .C1(_03157_),
    .C2(_03193_),
    .ZN(_04076_));
 NAND2_X1 _29251_ (.A1(_02654_),
    .A2(_02831_),
    .ZN(_04077_));
 NAND4_X1 _29252_ (.A1(_03211_),
    .A2(_02747_),
    .A3(_03234_),
    .A4(_02667_),
    .ZN(_04078_));
 NAND4_X1 _29253_ (.A1(_03211_),
    .A2(_03246_),
    .A3(_02684_),
    .A4(_03234_),
    .ZN(_04079_));
 NAND4_X1 _29254_ (.A1(_04077_),
    .A2(_03601_),
    .A3(_04078_),
    .A4(_04079_),
    .ZN(_04081_));
 AND4_X1 _29255_ (.A1(_03211_),
    .A2(_03148_),
    .A3(_03549_),
    .A4(_03234_),
    .ZN(_04082_));
 AOI211_X1 _29256_ (.A(_03149_),
    .B(_03189_),
    .C1(_02829_),
    .C2(_02657_),
    .ZN(_04083_));
 NOR4_X1 _29257_ (.A1(_04076_),
    .A2(_04081_),
    .A3(_04082_),
    .A4(_04083_),
    .ZN(_04084_));
 NAND4_X1 _29258_ (.A1(_04055_),
    .A2(_04066_),
    .A3(_04071_),
    .A4(_04084_),
    .ZN(_04085_));
 OAI21_X1 _29259_ (.A(_03541_),
    .B1(_03230_),
    .B2(_02658_),
    .ZN(_04086_));
 AND2_X1 _29260_ (.A1(_02765_),
    .A2(_02679_),
    .ZN(_04087_));
 AOI221_X4 _29261_ (.A(_04087_),
    .B1(_02796_),
    .B2(_02680_),
    .C1(_03528_),
    .C2(_03532_),
    .ZN(_04088_));
 OAI21_X1 _29262_ (.A(_03175_),
    .B1(_03160_),
    .B2(_02647_),
    .ZN(_04089_));
 AOI22_X1 _29263_ (.A1(_02703_),
    .A2(_03148_),
    .B1(_02765_),
    .B2(_03541_),
    .ZN(_04090_));
 AND4_X1 _29264_ (.A1(_04086_),
    .A2(_04088_),
    .A3(_04089_),
    .A4(_04090_),
    .ZN(_04091_));
 AND2_X1 _29265_ (.A1(_02629_),
    .A2(_02636_),
    .ZN(_04092_));
 OAI21_X1 _29266_ (.A(_02635_),
    .B1(_02641_),
    .B2(_04092_),
    .ZN(_04093_));
 OAI211_X1 _29267_ (.A(_04093_),
    .B(_03953_),
    .C1(_03155_),
    .C2(_03950_),
    .ZN(_04094_));
 OAI21_X1 _29268_ (.A(_02665_),
    .B1(_02641_),
    .B2(_02671_),
    .ZN(_04095_));
 NAND2_X1 _29269_ (.A1(_02665_),
    .A2(_03203_),
    .ZN(_04096_));
 NAND2_X1 _29270_ (.A1(_04095_),
    .A2(_04096_),
    .ZN(_04097_));
 NOR4_X1 _29271_ (.A1(_04094_),
    .A2(_04097_),
    .A3(_03580_),
    .A4(_03943_),
    .ZN(_04098_));
 NAND2_X1 _29272_ (.A1(_02717_),
    .A2(_02800_),
    .ZN(_04099_));
 OAI211_X1 _29273_ (.A(_02722_),
    .B(_02667_),
    .C1(_02829_),
    .C2(_02642_),
    .ZN(_04100_));
 OAI21_X1 _29274_ (.A(_02723_),
    .B1(_02670_),
    .B2(_02734_),
    .ZN(_04101_));
 AND3_X1 _29275_ (.A1(_04100_),
    .A2(_03575_),
    .A3(_04101_),
    .ZN(_04102_));
 OAI21_X1 _29276_ (.A(_02717_),
    .B1(_02727_),
    .B2(_02813_),
    .ZN(_04103_));
 OAI21_X1 _29277_ (.A(_02717_),
    .B1(_03209_),
    .B2(_03952_),
    .ZN(_04104_));
 AND4_X1 _29278_ (.A1(_04099_),
    .A2(_04102_),
    .A3(_04103_),
    .A4(_04104_),
    .ZN(_04105_));
 NAND2_X1 _29279_ (.A1(_02765_),
    .A2(_02731_),
    .ZN(_04106_));
 OAI21_X1 _29280_ (.A(_02742_),
    .B1(_02724_),
    .B2(_03209_),
    .ZN(_04107_));
 OAI21_X1 _29281_ (.A(_02733_),
    .B1(_02686_),
    .B2(_02654_),
    .ZN(_04108_));
 NAND2_X1 _29282_ (.A1(_02641_),
    .A2(_02736_),
    .ZN(_04109_));
 AND4_X1 _29283_ (.A1(_04106_),
    .A2(_04107_),
    .A3(_04108_),
    .A4(_04109_),
    .ZN(_04110_));
 NAND4_X1 _29284_ (.A1(_04091_),
    .A2(_04098_),
    .A3(_04105_),
    .A4(_04110_),
    .ZN(_04111_));
 NOR2_X2 _29285_ (.A1(_04085_),
    .A2(_04111_),
    .ZN(_04112_));
 XNOR2_X1 _29286_ (.A(_04112_),
    .B(_02837_),
    .ZN(_04113_));
 AND2_X1 _29287_ (.A1(_02534_),
    .A2(_02926_),
    .ZN(_04114_));
 AOI21_X1 _29288_ (.A(_03822_),
    .B1(_02444_),
    .B2(_02490_),
    .ZN(_04115_));
 AOI211_X1 _29289_ (.A(_04114_),
    .B(_04115_),
    .C1(_02468_),
    .C2(_02534_),
    .ZN(_04116_));
 OAI21_X1 _29290_ (.A(_02561_),
    .B1(_02563_),
    .B2(_02468_),
    .ZN(_04117_));
 AND4_X1 _29291_ (.A1(_02949_),
    .A2(_04116_),
    .A3(_02951_),
    .A4(_04117_),
    .ZN(_04118_));
 AOI21_X1 _29292_ (.A(_02938_),
    .B1(_03293_),
    .B2(_02409_),
    .ZN(_04119_));
 AOI21_X1 _29293_ (.A(_04119_),
    .B1(_02406_),
    .B2(_02549_),
    .ZN(_04120_));
 AOI211_X1 _29294_ (.A(_02956_),
    .B(_03839_),
    .C1(_02404_),
    .C2(_02540_),
    .ZN(_04122_));
 AND4_X1 _29295_ (.A1(_02539_),
    .A2(_04120_),
    .A3(_02542_),
    .A4(_04122_),
    .ZN(_04123_));
 OAI21_X1 _29296_ (.A(_02462_),
    .B1(_02541_),
    .B2(_02523_),
    .ZN(_04124_));
 AND3_X1 _29297_ (.A1(_04124_),
    .A2(_02463_),
    .A3(_03849_),
    .ZN(_04125_));
 OAI21_X1 _29298_ (.A(_02442_),
    .B1(_02609_),
    .B2(_02495_),
    .ZN(_04126_));
 AND4_X1 _29299_ (.A1(_02456_),
    .A2(_04125_),
    .A3(_02874_),
    .A4(_04126_),
    .ZN(_04127_));
 NAND4_X1 _29300_ (.A1(_03295_),
    .A2(_02397_),
    .A3(_02435_),
    .A4(_02438_),
    .ZN(_04128_));
 OAI211_X1 _29301_ (.A(_03292_),
    .B(_04128_),
    .C1(_02885_),
    .C2(_02933_),
    .ZN(_04129_));
 NAND4_X1 _29302_ (.A1(_03322_),
    .A2(_02557_),
    .A3(_02438_),
    .A4(_02558_),
    .ZN(_04130_));
 OAI21_X1 _29303_ (.A(_04130_),
    .B1(_02419_),
    .B2(_02572_),
    .ZN(_04131_));
 NAND3_X1 _29304_ (.A1(_02489_),
    .A2(_02586_),
    .A3(_02438_),
    .ZN(_04133_));
 NAND3_X1 _29305_ (.A1(_02404_),
    .A2(_02586_),
    .A3(_02389_),
    .ZN(_04134_));
 OAI211_X1 _29306_ (.A(_04133_),
    .B(_04134_),
    .C1(_02885_),
    .C2(_02572_),
    .ZN(_04135_));
 NOR4_X1 _29307_ (.A1(_04129_),
    .A2(_03303_),
    .A3(_04131_),
    .A4(_04135_),
    .ZN(_04136_));
 NAND4_X1 _29308_ (.A1(_04118_),
    .A2(_04123_),
    .A3(_04127_),
    .A4(_04136_),
    .ZN(_04137_));
 AOI21_X1 _29309_ (.A(_02569_),
    .B1(_02490_),
    .B2(_02544_),
    .ZN(_04138_));
 AOI21_X1 _29310_ (.A(_04138_),
    .B1(_02581_),
    .B2(_02578_),
    .ZN(_04139_));
 AND2_X1 _29311_ (.A1(_02575_),
    .A2(_02398_),
    .ZN(_04140_));
 INV_X1 _29312_ (.A(_04140_),
    .ZN(_04141_));
 AND3_X1 _29313_ (.A1(_04141_),
    .A2(_02576_),
    .A3(_02577_),
    .ZN(_04142_));
 OAI21_X1 _29314_ (.A(_02575_),
    .B1(_02410_),
    .B2(_02468_),
    .ZN(_04144_));
 AND4_X1 _29315_ (.A1(_02914_),
    .A2(_04139_),
    .A3(_04142_),
    .A4(_04144_),
    .ZN(_04145_));
 OAI21_X1 _29316_ (.A(_02600_),
    .B1(_02448_),
    .B2(_02489_),
    .ZN(_04146_));
 NAND2_X1 _29317_ (.A1(_02600_),
    .A2(_02564_),
    .ZN(_04147_));
 NAND3_X1 _29318_ (.A1(_02541_),
    .A2(_02437_),
    .A3(_02596_),
    .ZN(_04148_));
 NAND4_X1 _29319_ (.A1(_04146_),
    .A2(_02604_),
    .A3(_04147_),
    .A4(_04148_),
    .ZN(_04149_));
 AND2_X1 _29320_ (.A1(_02593_),
    .A2(_02465_),
    .ZN(_04150_));
 AND2_X1 _29321_ (.A1(_02592_),
    .A2(_02887_),
    .ZN(_04151_));
 OR2_X1 _29322_ (.A1(_04150_),
    .A2(_04151_),
    .ZN(_04152_));
 NAND4_X1 _29323_ (.A1(_02596_),
    .A2(_02880_),
    .A3(_02454_),
    .A4(_02554_),
    .ZN(_04153_));
 OAI21_X1 _29324_ (.A(_04153_),
    .B1(_02612_),
    .B2(_03832_),
    .ZN(_04155_));
 NAND2_X1 _29325_ (.A1(_02593_),
    .A2(_02500_),
    .ZN(_04156_));
 NAND4_X1 _29326_ (.A1(_02596_),
    .A2(_02470_),
    .A3(_02452_),
    .A4(_02554_),
    .ZN(_04157_));
 OAI211_X1 _29327_ (.A(_04156_),
    .B(_04157_),
    .C1(_02612_),
    .C2(_03305_),
    .ZN(_04158_));
 NOR4_X1 _29328_ (.A1(_04149_),
    .A2(_04152_),
    .A3(_04155_),
    .A4(_04158_),
    .ZN(_04159_));
 NAND2_X1 _29329_ (.A1(_02504_),
    .A2(_02578_),
    .ZN(_04160_));
 OAI211_X1 _29330_ (.A(_03865_),
    .B(_04160_),
    .C1(_03363_),
    .C2(_03894_),
    .ZN(_04161_));
 NAND3_X1 _29331_ (.A1(_02420_),
    .A2(_03295_),
    .A3(_02524_),
    .ZN(_04162_));
 OAI211_X1 _29332_ (.A(_04162_),
    .B(_03867_),
    .C1(_03363_),
    .C2(_02411_),
    .ZN(_04163_));
 NAND2_X1 _29333_ (.A1(_02483_),
    .A2(_02498_),
    .ZN(_04164_));
 INV_X1 _29334_ (.A(_02926_),
    .ZN(_04166_));
 OAI21_X1 _29335_ (.A(_04164_),
    .B1(_04166_),
    .B2(_03368_),
    .ZN(_04167_));
 OAI21_X1 _29336_ (.A(_03366_),
    .B1(_02544_),
    .B2(_03368_),
    .ZN(_04168_));
 NOR4_X1 _29337_ (.A1(_04161_),
    .A2(_04163_),
    .A3(_04167_),
    .A4(_04168_),
    .ZN(_04169_));
 NOR2_X1 _29338_ (.A1(_02485_),
    .A2(_02423_),
    .ZN(_04170_));
 AND2_X1 _29339_ (.A1(_02514_),
    .A2(_04170_),
    .ZN(_04171_));
 INV_X1 _29340_ (.A(_04171_),
    .ZN(_04172_));
 NAND3_X1 _29341_ (.A1(_02605_),
    .A2(_02927_),
    .A3(_02515_),
    .ZN(_04173_));
 NAND2_X1 _29342_ (.A1(_02515_),
    .A2(_02541_),
    .ZN(_04174_));
 AND3_X1 _29343_ (.A1(_04173_),
    .A2(_02525_),
    .A3(_04174_),
    .ZN(_04175_));
 NAND2_X1 _29344_ (.A1(_02905_),
    .A2(_02515_),
    .ZN(_04177_));
 OAI211_X1 _29345_ (.A(_02479_),
    .B(_03322_),
    .C1(_02880_),
    .C2(_02430_),
    .ZN(_04178_));
 NAND2_X1 _29346_ (.A1(_02479_),
    .A2(_02523_),
    .ZN(_04179_));
 NAND4_X1 _29347_ (.A1(_02397_),
    .A2(_02435_),
    .A3(_02524_),
    .A4(_02554_),
    .ZN(_04180_));
 AND3_X1 _29348_ (.A1(_04178_),
    .A2(_04179_),
    .A3(_04180_),
    .ZN(_04181_));
 AND4_X1 _29349_ (.A1(_04172_),
    .A2(_04175_),
    .A3(_04177_),
    .A4(_04181_),
    .ZN(_04182_));
 NAND4_X1 _29350_ (.A1(_04145_),
    .A2(_04159_),
    .A3(_04169_),
    .A4(_04182_),
    .ZN(_04183_));
 NOR2_X2 _29351_ (.A1(_04137_),
    .A2(_04183_),
    .ZN(_04184_));
 AOI21_X1 _29352_ (.A(_02125_),
    .B1(_02078_),
    .B2(_02020_),
    .ZN(_04185_));
 OAI21_X1 _29353_ (.A(_03800_),
    .B1(_02125_),
    .B2(_02107_),
    .ZN(_04186_));
 AND2_X1 _29354_ (.A1(_01952_),
    .A2(_01858_),
    .ZN(_04188_));
 AND3_X1 _29355_ (.A1(_01968_),
    .A2(_03003_),
    .A3(_01932_),
    .ZN(_04189_));
 NOR4_X1 _29356_ (.A1(_04185_),
    .A2(_04186_),
    .A3(_04188_),
    .A4(_04189_),
    .ZN(_04190_));
 NAND3_X1 _29357_ (.A1(_01992_),
    .A2(_01922_),
    .A3(_01852_),
    .ZN(_04191_));
 AND4_X1 _29358_ (.A1(_02061_),
    .A2(_01856_),
    .A3(_01932_),
    .A4(_01875_),
    .ZN(_04192_));
 AND2_X1 _29359_ (.A1(_02001_),
    .A2(_01992_),
    .ZN(_04193_));
 AOI211_X1 _29360_ (.A(_04192_),
    .B(_04193_),
    .C1(_01903_),
    .C2(_01992_),
    .ZN(_04194_));
 AND4_X1 _29361_ (.A1(_03430_),
    .A2(_04190_),
    .A3(_04191_),
    .A4(_04194_),
    .ZN(_04195_));
 AND4_X1 _29362_ (.A1(_01885_),
    .A2(_01922_),
    .A3(_02103_),
    .A4(_01887_),
    .ZN(_04196_));
 AND2_X1 _29363_ (.A1(_01890_),
    .A2(_01956_),
    .ZN(_04197_));
 AOI211_X1 _29364_ (.A(_04196_),
    .B(_04197_),
    .C1(_01890_),
    .C2(_01949_),
    .ZN(_04199_));
 OAI211_X1 _29365_ (.A(_03002_),
    .B(_01887_),
    .C1(_03401_),
    .C2(_01903_),
    .ZN(_04200_));
 OAI21_X1 _29366_ (.A(_01843_),
    .B1(_01911_),
    .B2(_01903_),
    .ZN(_04201_));
 NAND2_X1 _29367_ (.A1(_01843_),
    .A2(_02000_),
    .ZN(_04202_));
 NAND4_X1 _29368_ (.A1(_01928_),
    .A2(_03002_),
    .A3(_01995_),
    .A4(_01841_),
    .ZN(_04203_));
 AND4_X1 _29369_ (.A1(_03787_),
    .A2(_04201_),
    .A3(_04202_),
    .A4(_04203_),
    .ZN(_04204_));
 AND4_X1 _29370_ (.A1(_02114_),
    .A2(_04199_),
    .A3(_04200_),
    .A4(_04204_),
    .ZN(_04205_));
 NAND2_X1 _29371_ (.A1(_02014_),
    .A2(_02032_),
    .ZN(_04206_));
 AND3_X1 _29372_ (.A1(_04206_),
    .A2(_02015_),
    .A3(_01863_),
    .ZN(_04207_));
 OAI21_X1 _29373_ (.A(_02992_),
    .B1(_02009_),
    .B2(_01927_),
    .ZN(_04208_));
 NAND2_X1 _29374_ (.A1(_04208_),
    .A2(_02047_),
    .ZN(_04210_));
 OAI21_X1 _29375_ (.A(_02014_),
    .B1(_02035_),
    .B2(_01911_),
    .ZN(_04211_));
 AND4_X1 _29376_ (.A1(_03017_),
    .A2(_04207_),
    .A3(_04210_),
    .A4(_04211_),
    .ZN(_04212_));
 OAI21_X1 _29377_ (.A(_01934_),
    .B1(_01996_),
    .B2(_02061_),
    .ZN(_04213_));
 OAI211_X1 _29378_ (.A(_02132_),
    .B(_01852_),
    .C1(_02088_),
    .C2(_03405_),
    .ZN(_04214_));
 OAI21_X1 _29379_ (.A(_02132_),
    .B1(_01968_),
    .B2(_03401_),
    .ZN(_04215_));
 OAI211_X1 _29380_ (.A(_01934_),
    .B(_02009_),
    .C1(_02103_),
    .C2(_01852_),
    .ZN(_04216_));
 AND4_X1 _29381_ (.A1(_04213_),
    .A2(_04214_),
    .A3(_04215_),
    .A4(_04216_),
    .ZN(_04217_));
 NAND4_X1 _29382_ (.A1(_04195_),
    .A2(_04205_),
    .A3(_04212_),
    .A4(_04217_),
    .ZN(_04218_));
 AND2_X1 _29383_ (.A1(_01973_),
    .A2(_02108_),
    .ZN(_04219_));
 AND2_X1 _29384_ (.A1(_01973_),
    .A2(_02033_),
    .ZN(_04221_));
 AOI211_X1 _29385_ (.A(_04219_),
    .B(_04221_),
    .C1(_02098_),
    .C2(_01973_),
    .ZN(_04222_));
 OAI21_X1 _29386_ (.A(_01983_),
    .B1(_02076_),
    .B2(_02042_),
    .ZN(_04223_));
 OAI21_X1 _29387_ (.A(_01983_),
    .B1(_02032_),
    .B2(_02033_),
    .ZN(_04224_));
 AND4_X1 _29388_ (.A1(_01909_),
    .A2(_04222_),
    .A3(_04223_),
    .A4(_04224_),
    .ZN(_04225_));
 NAND2_X1 _29389_ (.A1(_01873_),
    .A2(_03397_),
    .ZN(_04226_));
 OAI21_X1 _29390_ (.A(_03395_),
    .B1(_01884_),
    .B2(_02007_),
    .ZN(_04227_));
 OAI21_X1 _29391_ (.A(_03397_),
    .B1(_01968_),
    .B2(_02061_),
    .ZN(_04228_));
 OAI21_X1 _29392_ (.A(_03395_),
    .B1(_02037_),
    .B2(_02039_),
    .ZN(_04229_));
 AND4_X1 _29393_ (.A1(_04226_),
    .A2(_04227_),
    .A3(_04228_),
    .A4(_04229_),
    .ZN(_04230_));
 OAI21_X1 _29394_ (.A(_02031_),
    .B1(_01968_),
    .B2(_02035_),
    .ZN(_04232_));
 OAI21_X1 _29395_ (.A(_04232_),
    .B1(_03023_),
    .B2(_02101_),
    .ZN(_04233_));
 NAND2_X1 _29396_ (.A1(_02031_),
    .A2(_02012_),
    .ZN(_04234_));
 NAND3_X1 _29397_ (.A1(_02033_),
    .A2(_03003_),
    .A3(_03020_),
    .ZN(_04235_));
 OAI211_X1 _29398_ (.A(_04234_),
    .B(_04235_),
    .C1(_03023_),
    .C2(_03426_),
    .ZN(_04236_));
 AOI21_X1 _29399_ (.A(_01971_),
    .B1(_02992_),
    .B2(_01877_),
    .ZN(_04237_));
 NOR4_X1 _29400_ (.A1(_04233_),
    .A2(_04236_),
    .A3(_03408_),
    .A4(_04237_),
    .ZN(_04238_));
 AND2_X1 _29401_ (.A1(_01899_),
    .A2(_02975_),
    .ZN(_04239_));
 AND4_X1 _29402_ (.A1(_01954_),
    .A2(_01896_),
    .A3(_01938_),
    .A4(_01875_),
    .ZN(_04240_));
 AND4_X1 _29403_ (.A1(_02061_),
    .A2(_01907_),
    .A3(_01980_),
    .A4(_01875_),
    .ZN(_04241_));
 AOI211_X1 _29404_ (.A(_04240_),
    .B(_04241_),
    .C1(_02035_),
    .C2(_01898_),
    .ZN(_04243_));
 OAI21_X1 _29405_ (.A(_01961_),
    .B1(_02000_),
    .B2(_01858_),
    .ZN(_04244_));
 OAI21_X1 _29406_ (.A(_01961_),
    .B1(_02057_),
    .B2(_02035_),
    .ZN(_04245_));
 AND4_X1 _29407_ (.A1(_04239_),
    .A2(_04243_),
    .A3(_04244_),
    .A4(_04245_),
    .ZN(_04246_));
 NAND4_X1 _29408_ (.A1(_04225_),
    .A2(_04230_),
    .A3(_04238_),
    .A4(_04246_),
    .ZN(_04247_));
 NOR2_X2 _29409_ (.A1(_04218_),
    .A2(_04247_),
    .ZN(_04248_));
 XNOR2_X1 _29410_ (.A(_04184_),
    .B(_04248_),
    .ZN(_04249_));
 XNOR2_X1 _29411_ (.A(_04113_),
    .B(_04249_),
    .ZN(_04250_));
 XNOR2_X1 _29412_ (.A(_04047_),
    .B(_04250_),
    .ZN(_04251_));
 XOR2_X1 _29413_ (.A(_04251_),
    .B(_17157_),
    .Z(_04252_));
 MUX2_X1 _29414_ (.A(_03987_),
    .B(_04252_),
    .S(_01825_),
    .Z(_00712_));
 XOR2_X1 _29415_ (.A(_17158_),
    .B(_17028_),
    .Z(_04254_));
 AOI211_X1 _29416_ (.A(_03070_),
    .B(_03073_),
    .C1(_02176_),
    .C2(_02380_),
    .ZN(_04255_));
 NOR2_X1 _29417_ (.A1(_02355_),
    .A2(_03084_),
    .ZN(_04256_));
 INV_X1 _29418_ (.A(_04256_),
    .ZN(_04257_));
 AND2_X1 _29419_ (.A1(_02247_),
    .A2(_02180_),
    .ZN(_04258_));
 AND2_X1 _29420_ (.A1(_02193_),
    .A2(_02180_),
    .ZN(_04259_));
 AND2_X1 _29421_ (.A1(_02222_),
    .A2(_02180_),
    .ZN(_04260_));
 NOR4_X1 _29422_ (.A1(_04258_),
    .A2(_04259_),
    .A3(_04013_),
    .A4(_04260_),
    .ZN(_04261_));
 OAI21_X1 _29423_ (.A(_02292_),
    .B1(_02309_),
    .B2(_02225_),
    .ZN(_04262_));
 AND4_X1 _29424_ (.A1(_04257_),
    .A2(_04261_),
    .A3(_03518_),
    .A4(_04262_),
    .ZN(_04264_));
 OAI221_X1 _29425_ (.A(_02380_),
    .B1(_03075_),
    .B2(_03080_),
    .C1(_02275_),
    .C2(_02352_),
    .ZN(_04265_));
 NAND2_X1 _29426_ (.A1(_02326_),
    .A2(_02204_),
    .ZN(_04266_));
 OAI21_X1 _29427_ (.A(_02325_),
    .B1(_03699_),
    .B2(_02318_),
    .ZN(_04267_));
 NAND4_X1 _29428_ (.A1(_02146_),
    .A2(_02259_),
    .A3(_02179_),
    .A4(_02260_),
    .ZN(_04268_));
 AND4_X1 _29429_ (.A1(_04266_),
    .A2(_04267_),
    .A3(_03078_),
    .A4(_04268_),
    .ZN(_04269_));
 AND4_X1 _29430_ (.A1(_04255_),
    .A2(_04264_),
    .A3(_04265_),
    .A4(_04269_),
    .ZN(_04270_));
 AND2_X1 _29431_ (.A1(_02363_),
    .A2(_02220_),
    .ZN(_04271_));
 AOI221_X4 _29432_ (.A(_03485_),
    .B1(_02143_),
    .B2(_02230_),
    .C1(_02259_),
    .C2(_02239_),
    .ZN(_04272_));
 NAND3_X1 _29433_ (.A1(_02347_),
    .A2(_02226_),
    .A3(_02227_),
    .ZN(_04273_));
 NAND2_X1 _29434_ (.A1(_03057_),
    .A2(_04273_),
    .ZN(_04275_));
 OR4_X1 _29435_ (.A1(_04271_),
    .A2(_04272_),
    .A3(_04022_),
    .A4(_04275_),
    .ZN(_04276_));
 INV_X1 _29436_ (.A(_02199_),
    .ZN(_04277_));
 AOI21_X1 _29437_ (.A(_02299_),
    .B1(_04277_),
    .B2(_02357_),
    .ZN(_04278_));
 AND2_X1 _29438_ (.A1(_02204_),
    .A2(_02238_),
    .ZN(_04279_));
 AND2_X1 _29439_ (.A1(_02378_),
    .A2(_02238_),
    .ZN(_04280_));
 OR4_X1 _29440_ (.A1(_03050_),
    .A2(_04278_),
    .A3(_04279_),
    .A4(_04280_),
    .ZN(_04281_));
 AND2_X1 _29441_ (.A1(_03062_),
    .A2(_02330_),
    .ZN(_04282_));
 INV_X1 _29442_ (.A(_04282_),
    .ZN(_04283_));
 NAND3_X1 _29443_ (.A1(_02318_),
    .A2(_02150_),
    .A3(_02227_),
    .ZN(_04284_));
 NAND2_X1 _29444_ (.A1(_02365_),
    .A2(_02357_),
    .ZN(_04286_));
 OAI21_X1 _29445_ (.A(_02152_),
    .B1(_04286_),
    .B2(_02304_),
    .ZN(_04287_));
 OAI21_X1 _29446_ (.A(_02334_),
    .B1(_02268_),
    .B2(_02347_),
    .ZN(_04288_));
 NAND4_X1 _29447_ (.A1(_04283_),
    .A2(_04284_),
    .A3(_04287_),
    .A4(_04288_),
    .ZN(_04289_));
 OAI21_X1 _29448_ (.A(_03483_),
    .B1(_03095_),
    .B2(_02299_),
    .ZN(_04290_));
 NOR4_X1 _29449_ (.A1(_04276_),
    .A2(_04281_),
    .A3(_04289_),
    .A4(_04290_),
    .ZN(_04291_));
 AOI211_X1 _29450_ (.A(_02185_),
    .B(_03093_),
    .C1(_03075_),
    .C2(_02285_),
    .ZN(_04292_));
 AOI21_X1 _29451_ (.A(_03093_),
    .B1(_03462_),
    .B2(_02205_),
    .ZN(_04293_));
 NOR3_X1 _29452_ (.A1(_04292_),
    .A2(_03715_),
    .A3(_04293_),
    .ZN(_04294_));
 NAND2_X1 _29453_ (.A1(_02192_),
    .A2(_03056_),
    .ZN(_04295_));
 OAI21_X1 _29454_ (.A(_04295_),
    .B1(_03114_),
    .B2(_03458_),
    .ZN(_04297_));
 AOI21_X1 _29455_ (.A(_03114_),
    .B1(_02203_),
    .B2(_02250_),
    .ZN(_04298_));
 AOI211_X1 _29456_ (.A(_04297_),
    .B(_04298_),
    .C1(_02192_),
    .C2(_03703_),
    .ZN(_04299_));
 OAI21_X1 _29457_ (.A(_02369_),
    .B1(_02248_),
    .B2(_02336_),
    .ZN(_04300_));
 AND3_X1 _29458_ (.A1(_04300_),
    .A2(_02289_),
    .A3(_02286_),
    .ZN(_04301_));
 INV_X1 _29459_ (.A(_02321_),
    .ZN(_04302_));
 NAND2_X1 _29460_ (.A1(_02209_),
    .A2(_02276_),
    .ZN(_04303_));
 AND4_X1 _29461_ (.A1(_03719_),
    .A2(_03107_),
    .A3(_04302_),
    .A4(_04303_),
    .ZN(_04304_));
 AND4_X1 _29462_ (.A1(_04294_),
    .A2(_04299_),
    .A3(_04301_),
    .A4(_04304_),
    .ZN(_04305_));
 AOI211_X1 _29463_ (.A(_02302_),
    .B(_04037_),
    .C1(_02328_),
    .C2(_02265_),
    .ZN(_04306_));
 NAND2_X1 _29464_ (.A1(_02254_),
    .A2(_02308_),
    .ZN(_04308_));
 AOI211_X1 _29465_ (.A(_02307_),
    .B(_03126_),
    .C1(_02345_),
    .C2(_02274_),
    .ZN(_04309_));
 NAND2_X1 _29466_ (.A1(_02274_),
    .A2(_02309_),
    .ZN(_04310_));
 OAI21_X1 _29467_ (.A(_02233_),
    .B1(_02193_),
    .B2(_02195_),
    .ZN(_04311_));
 NAND2_X1 _29468_ (.A1(_02311_),
    .A2(_02234_),
    .ZN(_04312_));
 NAND2_X1 _29469_ (.A1(_02234_),
    .A2(_02294_),
    .ZN(_04313_));
 AND3_X1 _29470_ (.A1(_04311_),
    .A2(_04312_),
    .A3(_04313_),
    .ZN(_04314_));
 AND4_X1 _29471_ (.A1(_04308_),
    .A2(_04309_),
    .A3(_04310_),
    .A4(_04314_),
    .ZN(_04315_));
 AND2_X1 _29472_ (.A1(_02157_),
    .A2(_02301_),
    .ZN(_04316_));
 OAI21_X1 _29473_ (.A(_02265_),
    .B1(_02200_),
    .B2(_04316_),
    .ZN(_04317_));
 OAI211_X1 _29474_ (.A(_02260_),
    .B(_02261_),
    .C1(_02294_),
    .C2(_02361_),
    .ZN(_04319_));
 AND4_X1 _29475_ (.A1(_02253_),
    .A2(_04033_),
    .A3(_02256_),
    .A4(_04319_),
    .ZN(_04320_));
 AND4_X1 _29476_ (.A1(_04306_),
    .A2(_04315_),
    .A3(_04317_),
    .A4(_04320_),
    .ZN(_04321_));
 AND4_X1 _29477_ (.A1(_04270_),
    .A2(_04291_),
    .A3(_04305_),
    .A4(_04321_),
    .ZN(_04322_));
 NAND2_X2 _29478_ (.A1(_04322_),
    .A2(_02283_),
    .ZN(_04323_));
 XOR2_X1 _29479_ (.A(_04323_),
    .B(_04248_),
    .Z(_04324_));
 AND2_X1 _29480_ (.A1(_01926_),
    .A2(_01902_),
    .ZN(_04325_));
 AOI211_X1 _29481_ (.A(_01919_),
    .B(_03386_),
    .C1(_02088_),
    .C2(_03405_),
    .ZN(_04326_));
 AOI211_X1 _29482_ (.A(_04325_),
    .B(_04326_),
    .C1(_01911_),
    .C2(_01983_),
    .ZN(_04327_));
 AND4_X1 _29483_ (.A1(_01894_),
    .A2(_01851_),
    .A3(_01980_),
    .A4(_01841_),
    .ZN(_04328_));
 AOI211_X1 _29484_ (.A(_04328_),
    .B(_04221_),
    .C1(_01973_),
    .C2(_02012_),
    .ZN(_04330_));
 OAI21_X1 _29485_ (.A(_01973_),
    .B1(_02035_),
    .B2(_03401_),
    .ZN(_04331_));
 OAI21_X1 _29486_ (.A(_01983_),
    .B1(_02098_),
    .B2(_01928_),
    .ZN(_04332_));
 NAND4_X1 _29487_ (.A1(_04327_),
    .A2(_04330_),
    .A3(_04331_),
    .A4(_04332_),
    .ZN(_04333_));
 OAI21_X1 _29488_ (.A(_01898_),
    .B1(_02079_),
    .B2(_02006_),
    .ZN(_04334_));
 NAND2_X1 _29489_ (.A1(_02076_),
    .A2(_01961_),
    .ZN(_04335_));
 NAND2_X1 _29490_ (.A1(_01898_),
    .A2(_01858_),
    .ZN(_04336_));
 OAI21_X1 _29491_ (.A(_01961_),
    .B1(_01949_),
    .B2(_01945_),
    .ZN(_04337_));
 NAND4_X1 _29492_ (.A1(_04334_),
    .A2(_04335_),
    .A3(_04336_),
    .A4(_04337_),
    .ZN(_04338_));
 NAND3_X1 _29493_ (.A1(_02059_),
    .A2(_01935_),
    .A3(_02009_),
    .ZN(_04339_));
 NAND2_X1 _29494_ (.A1(_02059_),
    .A2(_01953_),
    .ZN(_04341_));
 OAI211_X1 _29495_ (.A(_04339_),
    .B(_04341_),
    .C1(_01877_),
    .C2(_01971_),
    .ZN(_04342_));
 INV_X1 _29496_ (.A(_02053_),
    .ZN(_04343_));
 OAI21_X1 _29497_ (.A(_04343_),
    .B1(_03023_),
    .B2(_03390_),
    .ZN(_04344_));
 INV_X1 _29498_ (.A(_03791_),
    .ZN(_04345_));
 OAI21_X1 _29499_ (.A(_03407_),
    .B1(_04345_),
    .B2(_01971_),
    .ZN(_04346_));
 OAI211_X1 _29500_ (.A(_04234_),
    .B(_03410_),
    .C1(_03023_),
    .C2(_03426_),
    .ZN(_04347_));
 OR4_X1 _29501_ (.A1(_04342_),
    .A2(_04344_),
    .A3(_04346_),
    .A4(_04347_),
    .ZN(_04348_));
 OAI21_X1 _29502_ (.A(_03395_),
    .B1(_01915_),
    .B2(_01911_),
    .ZN(_04349_));
 OAI21_X1 _29503_ (.A(_03395_),
    .B1(_01873_),
    .B2(_02012_),
    .ZN(_04350_));
 AND2_X1 _29504_ (.A1(_04349_),
    .A2(_04350_),
    .ZN(_04352_));
 NAND2_X1 _29505_ (.A1(_02108_),
    .A2(_03397_),
    .ZN(_04353_));
 OAI211_X1 _29506_ (.A(_02018_),
    .B(_01852_),
    .C1(_02088_),
    .C2(_03405_),
    .ZN(_04354_));
 OAI21_X1 _29507_ (.A(_03397_),
    .B1(_02113_),
    .B2(_01939_),
    .ZN(_04355_));
 NAND4_X1 _29508_ (.A1(_04352_),
    .A2(_04353_),
    .A3(_04354_),
    .A4(_04355_),
    .ZN(_04356_));
 NOR4_X1 _29509_ (.A1(_04333_),
    .A2(_04338_),
    .A3(_04348_),
    .A4(_04356_),
    .ZN(_04357_));
 OAI22_X1 _29510_ (.A1(_02127_),
    .A2(_03405_),
    .B1(_02125_),
    .B2(_01990_),
    .ZN(_04358_));
 NOR2_X1 _29511_ (.A1(_01986_),
    .A2(_02125_),
    .ZN(_04359_));
 NOR4_X1 _29512_ (.A1(_02123_),
    .A2(_04358_),
    .A3(_04359_),
    .A4(_04188_),
    .ZN(_04360_));
 OAI221_X1 _29513_ (.A(_01992_),
    .B1(_01954_),
    .B2(_01920_),
    .C1(_02061_),
    .C2(_01905_),
    .ZN(_04361_));
 AND4_X1 _29514_ (.A1(_03430_),
    .A2(_04360_),
    .A3(_02987_),
    .A4(_04361_),
    .ZN(_04363_));
 NAND3_X1 _29515_ (.A1(_02132_),
    .A2(_01894_),
    .A3(_02103_),
    .ZN(_04364_));
 NAND2_X1 _29516_ (.A1(_02132_),
    .A2(_03401_),
    .ZN(_04365_));
 NAND4_X1 _29517_ (.A1(_02996_),
    .A2(_04364_),
    .A3(_01998_),
    .A4(_04365_),
    .ZN(_04366_));
 AOI21_X1 _29518_ (.A(_03439_),
    .B1(_03811_),
    .B2(_01919_),
    .ZN(_04367_));
 AND2_X1 _29519_ (.A1(_02986_),
    .A2(_01934_),
    .ZN(_04368_));
 NOR4_X1 _29520_ (.A1(_04366_),
    .A2(_04367_),
    .A3(_04368_),
    .A4(_03443_),
    .ZN(_04369_));
 AND4_X1 _29521_ (.A1(_03405_),
    .A2(_03002_),
    .A3(_01852_),
    .A4(_01875_),
    .ZN(_04370_));
 AND4_X1 _29522_ (.A1(_03002_),
    .A2(_01894_),
    .A3(_02103_),
    .A4(_01875_),
    .ZN(_04371_));
 AOI211_X1 _29523_ (.A(_04370_),
    .B(_04371_),
    .C1(_02046_),
    .C2(_02047_),
    .ZN(_04372_));
 NAND2_X1 _29524_ (.A1(_01890_),
    .A2(_02037_),
    .ZN(_04374_));
 OAI21_X1 _29525_ (.A(_01890_),
    .B1(_02108_),
    .B2(_01956_),
    .ZN(_04375_));
 AND4_X1 _29526_ (.A1(_04374_),
    .A2(_01913_),
    .A3(_04375_),
    .A4(_01916_),
    .ZN(_04376_));
 OAI21_X1 _29527_ (.A(_02014_),
    .B1(_02000_),
    .B2(_01949_),
    .ZN(_04377_));
 NAND4_X1 _29528_ (.A1(_03002_),
    .A2(_03003_),
    .A3(_01905_),
    .A4(_01922_),
    .ZN(_04378_));
 AND4_X1 _29529_ (.A1(_01859_),
    .A2(_04377_),
    .A3(_03808_),
    .A4(_04378_),
    .ZN(_04379_));
 NAND3_X1 _29530_ (.A1(_02039_),
    .A2(_03002_),
    .A3(_01841_),
    .ZN(_04380_));
 AND4_X1 _29531_ (.A1(_03010_),
    .A2(_03787_),
    .A3(_04202_),
    .A4(_04380_),
    .ZN(_04381_));
 AND4_X1 _29532_ (.A1(_04372_),
    .A2(_04376_),
    .A3(_04379_),
    .A4(_04381_),
    .ZN(_04382_));
 NAND4_X1 _29533_ (.A1(_04357_),
    .A2(_04363_),
    .A3(_04369_),
    .A4(_04382_),
    .ZN(_04383_));
 NOR2_X2 _29534_ (.A1(_04383_),
    .A2(_02045_),
    .ZN(_04385_));
 NAND4_X1 _29535_ (.A1(_02596_),
    .A2(_02470_),
    .A3(_02472_),
    .A4(_02558_),
    .ZN(_04386_));
 OAI21_X1 _29536_ (.A(_04386_),
    .B1(_02569_),
    .B2(_03823_),
    .ZN(_04387_));
 INV_X1 _29537_ (.A(_02482_),
    .ZN(_04388_));
 NAND2_X1 _29538_ (.A1(_02595_),
    .A2(_02479_),
    .ZN(_04389_));
 NAND3_X1 _29539_ (.A1(_04388_),
    .A2(_04389_),
    .A3(_04179_),
    .ZN(_04390_));
 AND4_X1 _29540_ (.A1(_02470_),
    .A2(_02472_),
    .A3(_02524_),
    .A4(_02554_),
    .ZN(_04391_));
 NAND2_X1 _29541_ (.A1(_02410_),
    .A2(_02549_),
    .ZN(_04392_));
 NAND2_X1 _29542_ (.A1(_02467_),
    .A2(_02549_),
    .ZN(_04393_));
 NAND2_X1 _29543_ (.A1(_04392_),
    .A2(_04393_),
    .ZN(_04394_));
 OR4_X1 _29544_ (.A1(_04387_),
    .A2(_04390_),
    .A3(_04391_),
    .A4(_04394_),
    .ZN(_04396_));
 AND2_X1 _29545_ (.A1(_02905_),
    .A2(_02514_),
    .ZN(_04397_));
 AND2_X1 _29546_ (.A1(_02514_),
    .A2(_03335_),
    .ZN(_04398_));
 OR4_X1 _29547_ (.A1(_02907_),
    .A2(_04397_),
    .A3(_02931_),
    .A4(_04398_),
    .ZN(_04399_));
 AOI21_X1 _29548_ (.A(_02516_),
    .B1(_03883_),
    .B2(_02414_),
    .ZN(_04400_));
 NOR4_X1 _29549_ (.A1(_04396_),
    .A2(_04399_),
    .A3(_02616_),
    .A4(_04400_),
    .ZN(_04401_));
 AOI211_X1 _29550_ (.A(_02414_),
    .B(_02588_),
    .C1(_02880_),
    .C2(_02430_),
    .ZN(_04402_));
 OAI21_X1 _29551_ (.A(_02540_),
    .B1(_02404_),
    .B2(_02571_),
    .ZN(_04403_));
 OAI21_X1 _29552_ (.A(_02540_),
    .B1(_02468_),
    .B2(_02523_),
    .ZN(_04404_));
 NAND4_X1 _29553_ (.A1(_02472_),
    .A2(_03322_),
    .A3(_02437_),
    .A4(_02553_),
    .ZN(_04405_));
 NAND3_X1 _29554_ (.A1(_04403_),
    .A2(_04404_),
    .A3(_04405_),
    .ZN(_04407_));
 OAI211_X1 _29555_ (.A(_02561_),
    .B(_02435_),
    .C1(_02428_),
    .C2(_02430_),
    .ZN(_04408_));
 NAND3_X1 _29556_ (.A1(_02578_),
    .A2(_02553_),
    .A3(_02558_),
    .ZN(_04409_));
 OAI21_X1 _29557_ (.A(_02561_),
    .B1(_02476_),
    .B2(_02527_),
    .ZN(_04410_));
 NAND3_X1 _29558_ (.A1(_04408_),
    .A2(_04409_),
    .A3(_04410_),
    .ZN(_04411_));
 NAND3_X1 _29559_ (.A1(_02489_),
    .A2(_03295_),
    .A3(_02596_),
    .ZN(_04412_));
 OAI211_X1 _29560_ (.A(_02579_),
    .B(_04412_),
    .C1(_02588_),
    .C2(_03305_),
    .ZN(_04413_));
 NOR4_X1 _29561_ (.A1(_04402_),
    .A2(_04407_),
    .A3(_04411_),
    .A4(_04413_),
    .ZN(_04414_));
 OAI22_X1 _29562_ (.A1(_03293_),
    .A2(_03822_),
    .B1(_02885_),
    .B2(_02572_),
    .ZN(_04415_));
 OAI21_X1 _29563_ (.A(_02504_),
    .B1(_02483_),
    .B2(_02468_),
    .ZN(_04416_));
 OAI21_X1 _29564_ (.A(_04416_),
    .B1(_03325_),
    .B2(_03363_),
    .ZN(_04418_));
 NAND2_X1 _29565_ (.A1(_02461_),
    .A2(_03882_),
    .ZN(_04419_));
 NAND2_X1 _29566_ (.A1(_02549_),
    .A2(_02541_),
    .ZN(_04420_));
 NAND3_X1 _29567_ (.A1(_02455_),
    .A2(_02437_),
    .A3(_02596_),
    .ZN(_04421_));
 NAND4_X1 _29568_ (.A1(_04156_),
    .A2(_04419_),
    .A3(_04420_),
    .A4(_04421_),
    .ZN(_04422_));
 NOR4_X1 _29569_ (.A1(_04415_),
    .A2(_04418_),
    .A3(_02585_),
    .A4(_04422_),
    .ZN(_04423_));
 OAI211_X1 _29570_ (.A(_04160_),
    .B(_03366_),
    .C1(_03822_),
    .C2(_02447_),
    .ZN(_04424_));
 NOR4_X1 _29571_ (.A1(_04424_),
    .A2(_02598_),
    .A3(_02552_),
    .A4(_03872_),
    .ZN(_04425_));
 NAND4_X1 _29572_ (.A1(_04401_),
    .A2(_04414_),
    .A3(_04423_),
    .A4(_04425_),
    .ZN(_04426_));
 AOI22_X1 _29573_ (.A1(_02600_),
    .A2(_02489_),
    .B1(_02391_),
    .B2(_02595_),
    .ZN(_04427_));
 OAI211_X1 _29574_ (.A(_04427_),
    .B(_03302_),
    .C1(_03894_),
    .C2(_02938_),
    .ZN(_04429_));
 OAI21_X1 _29575_ (.A(_02483_),
    .B1(_02549_),
    .B2(_02498_),
    .ZN(_04430_));
 NAND2_X1 _29576_ (.A1(_02602_),
    .A2(_02462_),
    .ZN(_04431_));
 NAND4_X1 _29577_ (.A1(_04430_),
    .A2(_02945_),
    .A3(_02919_),
    .A4(_04431_),
    .ZN(_04432_));
 NOR4_X1 _29578_ (.A1(_04429_),
    .A2(_02910_),
    .A3(_04432_),
    .A4(_04150_),
    .ZN(_04433_));
 OR2_X1 _29579_ (.A1(_02509_),
    .A2(_03888_),
    .ZN(_04434_));
 OAI21_X1 _29580_ (.A(_02432_),
    .B1(_04434_),
    .B2(_02470_),
    .ZN(_04435_));
 AOI22_X1 _29581_ (.A1(_03895_),
    .A2(_02504_),
    .B1(_02564_),
    .B2(_02600_),
    .ZN(_04436_));
 OAI21_X1 _29582_ (.A(_02462_),
    .B1(_02547_),
    .B2(_02887_),
    .ZN(_04437_));
 NAND2_X1 _29583_ (.A1(_02490_),
    .A2(_03308_),
    .ZN(_04438_));
 OAI21_X1 _29584_ (.A(_02391_),
    .B1(_04438_),
    .B2(_02495_),
    .ZN(_04440_));
 OAI21_X1 _29585_ (.A(_02442_),
    .B1(_02458_),
    .B2(_02571_),
    .ZN(_04441_));
 OAI21_X1 _29586_ (.A(_02442_),
    .B1(_02410_),
    .B2(_02595_),
    .ZN(_04442_));
 AND4_X1 _29587_ (.A1(_04437_),
    .A2(_04440_),
    .A3(_04441_),
    .A4(_04442_),
    .ZN(_04443_));
 NAND4_X1 _29588_ (.A1(_04433_),
    .A2(_04435_),
    .A3(_04436_),
    .A4(_04443_),
    .ZN(_04444_));
 NOR2_X2 _29589_ (.A1(_04426_),
    .A2(_04444_),
    .ZN(_04445_));
 XNOR2_X2 _29590_ (.A(_04385_),
    .B(_04445_),
    .ZN(_04446_));
 XNOR2_X1 _29591_ (.A(_04324_),
    .B(_04446_),
    .ZN(_04447_));
 AOI21_X1 _29592_ (.A(_03200_),
    .B1(_02816_),
    .B2(_02715_),
    .ZN(_04448_));
 AND4_X1 _29593_ (.A1(_02642_),
    .A2(_03211_),
    .A3(_02694_),
    .A4(_02702_),
    .ZN(_04449_));
 AND4_X1 _29594_ (.A1(_02674_),
    .A2(_02803_),
    .A3(_02694_),
    .A4(_02652_),
    .ZN(_04451_));
 OR4_X1 _29595_ (.A1(_03916_),
    .A2(_04448_),
    .A3(_04449_),
    .A4(_04451_),
    .ZN(_04452_));
 AND2_X1 _29596_ (.A1(_02812_),
    .A2(_02727_),
    .ZN(_04453_));
 NOR4_X1 _29597_ (.A1(_04452_),
    .A2(_03241_),
    .A3(_03611_),
    .A4(_04453_),
    .ZN(_04454_));
 OAI21_X1 _29598_ (.A(_02831_),
    .B1(_02720_),
    .B2(_02641_),
    .ZN(_04455_));
 OAI21_X1 _29599_ (.A(_02831_),
    .B1(_02711_),
    .B2(_02698_),
    .ZN(_04456_));
 NOR2_X1 _29600_ (.A1(_03193_),
    .A2(_03201_),
    .ZN(_04457_));
 NOR2_X1 _29601_ (.A1(_04457_),
    .A2(_04073_),
    .ZN(_04458_));
 AND4_X1 _29602_ (.A1(_03226_),
    .A2(_04455_),
    .A3(_04456_),
    .A4(_04458_),
    .ZN(_04459_));
 OAI21_X1 _29603_ (.A(_03172_),
    .B1(_03169_),
    .B2(_03209_),
    .ZN(_04460_));
 OAI21_X1 _29604_ (.A(_03172_),
    .B1(_02813_),
    .B2(_02728_),
    .ZN(_04462_));
 OAI211_X1 _29605_ (.A(_02759_),
    .B(_16778_),
    .C1(_16777_),
    .C2(_02638_),
    .ZN(_04463_));
 AND4_X1 _29606_ (.A1(_03177_),
    .A2(_04460_),
    .A3(_04462_),
    .A4(_04463_),
    .ZN(_04464_));
 OAI211_X1 _29607_ (.A(_02781_),
    .B(_02783_),
    .C1(_03145_),
    .C2(_03206_),
    .ZN(_04465_));
 NAND2_X1 _29608_ (.A1(_02670_),
    .A2(_02799_),
    .ZN(_04466_));
 OAI211_X1 _29609_ (.A(_04466_),
    .B(_04049_),
    .C1(_03206_),
    .C2(_03152_),
    .ZN(_04467_));
 INV_X1 _29610_ (.A(_03544_),
    .ZN(_04468_));
 AOI21_X1 _29611_ (.A(_03190_),
    .B1(_04468_),
    .B2(_03145_),
    .ZN(_04469_));
 NOR4_X1 _29612_ (.A1(_03924_),
    .A2(_04465_),
    .A3(_04467_),
    .A4(_04469_),
    .ZN(_04470_));
 NAND4_X1 _29613_ (.A1(_04454_),
    .A2(_04459_),
    .A3(_04464_),
    .A4(_04470_),
    .ZN(_04471_));
 OAI21_X1 _29614_ (.A(_02665_),
    .B1(_02818_),
    .B2(_02782_),
    .ZN(_04473_));
 OAI211_X1 _29615_ (.A(_02664_),
    .B(_02800_),
    .C1(_02829_),
    .C2(_02657_),
    .ZN(_04474_));
 AND3_X1 _29616_ (.A1(_04473_),
    .A2(_04096_),
    .A3(_04474_),
    .ZN(_04475_));
 OAI211_X1 _29617_ (.A(_03234_),
    .B(_02622_),
    .C1(_02675_),
    .C2(_02671_),
    .ZN(_04476_));
 NAND3_X1 _29618_ (.A1(_02737_),
    .A2(_03234_),
    .A3(_02622_),
    .ZN(_04477_));
 AND3_X1 _29619_ (.A1(_02659_),
    .A2(_03192_),
    .A3(_04477_),
    .ZN(_04478_));
 AND4_X1 _29620_ (.A1(_02634_),
    .A2(_04475_),
    .A3(_04476_),
    .A4(_04478_),
    .ZN(_04479_));
 OAI211_X1 _29621_ (.A(_03142_),
    .B(_02712_),
    .C1(_03145_),
    .C2(_02713_),
    .ZN(_04480_));
 AOI21_X1 _29622_ (.A(_03146_),
    .B1(_02816_),
    .B2(_04468_),
    .ZN(_04481_));
 AOI21_X1 _29623_ (.A(_02713_),
    .B1(_03152_),
    .B2(_03572_),
    .ZN(_04482_));
 NOR4_X1 _29624_ (.A1(_04480_),
    .A2(_03577_),
    .A3(_04481_),
    .A4(_04482_),
    .ZN(_04484_));
 OAI21_X1 _29625_ (.A(_03541_),
    .B1(_02670_),
    .B2(_02734_),
    .ZN(_04485_));
 NAND3_X1 _29626_ (.A1(_02680_),
    .A2(_02684_),
    .A3(_03549_),
    .ZN(_04486_));
 NAND2_X1 _29627_ (.A1(_02704_),
    .A2(_02680_),
    .ZN(_04487_));
 AND3_X1 _29628_ (.A1(_04486_),
    .A2(_04487_),
    .A3(_02681_),
    .ZN(_04488_));
 OAI21_X1 _29629_ (.A(_03175_),
    .B1(_03169_),
    .B2(_02686_),
    .ZN(_04489_));
 OAI21_X1 _29630_ (.A(_03541_),
    .B1(_02833_),
    .B2(_03952_),
    .ZN(_04490_));
 AND4_X1 _29631_ (.A1(_04485_),
    .A2(_04488_),
    .A3(_04489_),
    .A4(_04490_),
    .ZN(_04491_));
 AOI21_X1 _29632_ (.A(_03535_),
    .B1(_03948_),
    .B2(_03149_),
    .ZN(_04492_));
 NAND2_X1 _29633_ (.A1(_02670_),
    .A2(_02733_),
    .ZN(_04493_));
 NAND3_X1 _29634_ (.A1(_02733_),
    .A2(_02832_),
    .A3(_03246_),
    .ZN(_04495_));
 NAND2_X1 _29635_ (.A1(_02732_),
    .A2(_02643_),
    .ZN(_04496_));
 NAND3_X1 _29636_ (.A1(_04493_),
    .A2(_04495_),
    .A3(_04496_),
    .ZN(_04497_));
 NOR4_X1 _29637_ (.A1(_03163_),
    .A2(_03537_),
    .A3(_04492_),
    .A4(_04497_),
    .ZN(_04498_));
 NAND4_X1 _29638_ (.A1(_04479_),
    .A2(_04484_),
    .A3(_04491_),
    .A4(_04498_),
    .ZN(_04499_));
 NOR2_X2 _29639_ (.A1(_04471_),
    .A2(_04499_),
    .ZN(_04500_));
 XNOR2_X1 _29640_ (.A(_04447_),
    .B(_04500_),
    .ZN(_04501_));
 XNOR2_X1 _29641_ (.A(_04501_),
    .B(_17158_),
    .ZN(_04502_));
 MUX2_X1 _29642_ (.A(_04254_),
    .B(_04502_),
    .S(_01825_),
    .Z(_00713_));
 XOR2_X1 _29643_ (.A(_17159_),
    .B(_17030_),
    .Z(_04503_));
 OAI21_X1 _29644_ (.A(_01952_),
    .B1(_01956_),
    .B2(_01949_),
    .ZN(_04505_));
 OAI21_X1 _29645_ (.A(_01952_),
    .B1(_01968_),
    .B2(_03401_),
    .ZN(_04506_));
 NAND3_X1 _29646_ (.A1(_04505_),
    .A2(_04506_),
    .A3(_03799_),
    .ZN(_04507_));
 AND2_X1 _29647_ (.A1(_01947_),
    .A2(_01897_),
    .ZN(_04508_));
 AND2_X1 _29648_ (.A1(_01942_),
    .A2(_01948_),
    .ZN(_04509_));
 NAND2_X1 _29649_ (.A1(_01897_),
    .A2(_01902_),
    .ZN(_04510_));
 NAND2_X1 _29650_ (.A1(_02084_),
    .A2(_04510_),
    .ZN(_04511_));
 OR4_X1 _29651_ (.A1(_04509_),
    .A2(_03762_),
    .A3(_02982_),
    .A4(_04511_),
    .ZN(_04512_));
 AOI21_X1 _29652_ (.A(_03439_),
    .B1(_02068_),
    .B2(_01990_),
    .ZN(_04513_));
 NAND2_X1 _29653_ (.A1(_01870_),
    .A2(_01975_),
    .ZN(_04514_));
 INV_X1 _29654_ (.A(_01890_),
    .ZN(_04516_));
 OAI21_X1 _29655_ (.A(_04514_),
    .B1(_04516_),
    .B2(_03389_),
    .ZN(_04517_));
 OR4_X1 _29656_ (.A1(_04508_),
    .A2(_04512_),
    .A3(_04513_),
    .A4(_04517_),
    .ZN(_04518_));
 AND2_X1 _29657_ (.A1(_01855_),
    .A2(_01884_),
    .ZN(_04519_));
 OR3_X1 _29658_ (.A1(_04519_),
    .A2(_03375_),
    .A3(_04325_),
    .ZN(_04520_));
 AOI22_X1 _29659_ (.A1(_01963_),
    .A2(_01901_),
    .B1(_01933_),
    .B2(_01902_),
    .ZN(_04521_));
 OAI21_X1 _29660_ (.A(_01958_),
    .B1(_01956_),
    .B2(_01948_),
    .ZN(_04522_));
 NAND3_X1 _29661_ (.A1(_01924_),
    .A2(_01838_),
    .A3(_01886_),
    .ZN(_04523_));
 NAND4_X1 _29662_ (.A1(_04521_),
    .A2(_03430_),
    .A3(_04522_),
    .A4(_04523_),
    .ZN(_04524_));
 NAND2_X1 _29663_ (.A1(_01889_),
    .A2(_02098_),
    .ZN(_04525_));
 AOI22_X1 _29664_ (.A1(_01943_),
    .A2(_02012_),
    .B1(_01974_),
    .B2(_01847_),
    .ZN(_04527_));
 NAND4_X1 _29665_ (.A1(_02052_),
    .A2(_04525_),
    .A3(_02087_),
    .A4(_04527_),
    .ZN(_04528_));
 OR4_X1 _29666_ (.A1(_03425_),
    .A2(_04520_),
    .A3(_04524_),
    .A4(_04528_),
    .ZN(_04529_));
 NOR4_X1 _29667_ (.A1(_01937_),
    .A2(_01858_),
    .A3(_02037_),
    .A4(_02012_),
    .ZN(_04530_));
 OAI22_X1 _29668_ (.A1(_04530_),
    .A2(_03386_),
    .B1(_01946_),
    .B2(_03431_),
    .ZN(_04531_));
 OR4_X1 _29669_ (.A1(_04507_),
    .A2(_04518_),
    .A3(_04529_),
    .A4(_04531_),
    .ZN(_04532_));
 AOI22_X1 _29670_ (.A1(_01961_),
    .A2(_01945_),
    .B1(_01979_),
    .B2(_02132_),
    .ZN(_04533_));
 NAND2_X1 _29671_ (.A1(_01915_),
    .A2(_03395_),
    .ZN(_04534_));
 OAI211_X1 _29672_ (.A(_04533_),
    .B(_04534_),
    .C1(_02078_),
    .C2(_01971_),
    .ZN(_04535_));
 NAND2_X1 _29673_ (.A1(_02005_),
    .A2(_02061_),
    .ZN(_04536_));
 NOR2_X1 _29674_ (.A1(_04516_),
    .A2(_04536_),
    .ZN(_04538_));
 OAI221_X1 _29675_ (.A(_02996_),
    .B1(_02977_),
    .B2(_02077_),
    .C1(_02109_),
    .C2(_03439_),
    .ZN(_04539_));
 OAI211_X1 _29676_ (.A(_01882_),
    .B(_01841_),
    .C1(_01885_),
    .C2(_01896_),
    .ZN(_04540_));
 NAND4_X1 _29677_ (.A1(_04540_),
    .A2(_03806_),
    .A3(_03007_),
    .A4(_03394_),
    .ZN(_04541_));
 OR4_X1 _29678_ (.A1(_04538_),
    .A2(_04539_),
    .A3(_04541_),
    .A4(_01864_),
    .ZN(_04542_));
 OAI21_X1 _29679_ (.A(_02059_),
    .B1(_02110_),
    .B2(_02113_),
    .ZN(_04543_));
 OAI211_X1 _29680_ (.A(_02018_),
    .B(_01852_),
    .C1(_01954_),
    .C2(_03405_),
    .ZN(_04544_));
 OAI21_X1 _29681_ (.A(_02018_),
    .B1(_02001_),
    .B2(_02042_),
    .ZN(_04545_));
 OAI21_X1 _29682_ (.A(_02992_),
    .B1(_01919_),
    .B2(_01846_),
    .ZN(_04546_));
 AOI22_X1 _29683_ (.A1(_04546_),
    .A2(_01898_),
    .B1(_01961_),
    .B2(_02057_),
    .ZN(_04547_));
 NAND4_X1 _29684_ (.A1(_04543_),
    .A2(_04544_),
    .A3(_04545_),
    .A4(_04547_),
    .ZN(_04549_));
 AOI21_X1 _29685_ (.A(_01879_),
    .B1(_03757_),
    .B2(_04345_),
    .ZN(_04550_));
 AOI21_X1 _29686_ (.A(_04550_),
    .B1(_01937_),
    .B2(_02047_),
    .ZN(_04551_));
 OAI21_X1 _29687_ (.A(_02031_),
    .B1(_02042_),
    .B2(_03791_),
    .ZN(_04552_));
 NAND4_X1 _29688_ (.A1(_01928_),
    .A2(_02094_),
    .A3(_01995_),
    .A4(_03020_),
    .ZN(_04553_));
 NAND4_X1 _29689_ (.A1(_02094_),
    .A2(_01851_),
    .A3(_01920_),
    .A4(_03020_),
    .ZN(_04554_));
 AND3_X1 _29690_ (.A1(_04552_),
    .A2(_04553_),
    .A3(_04554_),
    .ZN(_04555_));
 NAND2_X1 _29691_ (.A1(_01843_),
    .A2(_02012_),
    .ZN(_04556_));
 OAI22_X1 _29692_ (.A1(_01893_),
    .A2(_01954_),
    .B1(_02009_),
    .B2(_01927_),
    .ZN(_04557_));
 OAI21_X1 _29693_ (.A(_01843_),
    .B1(_04557_),
    .B2(_01979_),
    .ZN(_04558_));
 NAND4_X1 _29694_ (.A1(_04551_),
    .A2(_04555_),
    .A3(_04556_),
    .A4(_04558_),
    .ZN(_04560_));
 OR4_X1 _29695_ (.A1(_04535_),
    .A2(_04542_),
    .A3(_04549_),
    .A4(_04560_),
    .ZN(_04561_));
 NOR2_X2 _29696_ (.A1(_04532_),
    .A2(_04561_),
    .ZN(_04562_));
 AND4_X1 _29697_ (.A1(_02470_),
    .A2(_02553_),
    .A3(_02423_),
    .A4(_02554_),
    .ZN(_04563_));
 AND2_X1 _29698_ (.A1(_02548_),
    .A2(_02570_),
    .ZN(_04564_));
 AOI211_X1 _29699_ (.A(_04563_),
    .B(_04564_),
    .C1(_02509_),
    .C2(_02549_),
    .ZN(_04565_));
 OAI21_X1 _29700_ (.A(_02561_),
    .B1(_02448_),
    .B2(_02897_),
    .ZN(_04566_));
 AND3_X1 _29701_ (.A1(_02481_),
    .A2(_02532_),
    .A3(_02417_),
    .ZN(_04567_));
 AND2_X1 _29702_ (.A1(_02560_),
    .A2(_02476_),
    .ZN(_04568_));
 AOI211_X1 _29703_ (.A(_04567_),
    .B(_04568_),
    .C1(_02561_),
    .C2(_03888_),
    .ZN(_04569_));
 OAI211_X1 _29704_ (.A(_03295_),
    .B(_02553_),
    .C1(_02446_),
    .C2(_02495_),
    .ZN(_04571_));
 OAI21_X1 _29705_ (.A(_02534_),
    .B1(_02926_),
    .B2(_02466_),
    .ZN(_04572_));
 AND4_X1 _29706_ (.A1(_04566_),
    .A2(_04569_),
    .A3(_04571_),
    .A4(_04572_),
    .ZN(_04573_));
 OAI211_X1 _29707_ (.A(_02549_),
    .B(_16730_),
    .C1(_02880_),
    .C2(_02392_),
    .ZN(_04574_));
 NAND2_X1 _29708_ (.A1(_02540_),
    .A2(_02523_),
    .ZN(_04575_));
 NAND2_X1 _29709_ (.A1(_02540_),
    .A2(_02446_),
    .ZN(_04576_));
 AND4_X1 _29710_ (.A1(_02959_),
    .A2(_03840_),
    .A3(_04575_),
    .A4(_04576_),
    .ZN(_04577_));
 AND4_X1 _29711_ (.A1(_04565_),
    .A2(_04573_),
    .A3(_04574_),
    .A4(_04577_),
    .ZN(_04578_));
 OAI21_X1 _29712_ (.A(_02504_),
    .B1(_02500_),
    .B2(_02450_),
    .ZN(_04579_));
 OAI21_X1 _29713_ (.A(_02504_),
    .B1(_02420_),
    .B2(_02523_),
    .ZN(_04580_));
 AND3_X1 _29714_ (.A1(_04579_),
    .A2(_04580_),
    .A3(_03866_),
    .ZN(_04582_));
 AND2_X1 _29715_ (.A1(_02486_),
    .A2(_02493_),
    .ZN(_04583_));
 AOI211_X1 _29716_ (.A(_04583_),
    .B(_03360_),
    .C1(_03322_),
    .C2(_02498_),
    .ZN(_04584_));
 NAND2_X1 _29717_ (.A1(_02515_),
    .A2(_02468_),
    .ZN(_04585_));
 NAND2_X1 _29718_ (.A1(_02514_),
    .A2(_02500_),
    .ZN(_04586_));
 AND4_X1 _29719_ (.A1(_04585_),
    .A2(_04586_),
    .A3(_03898_),
    .A4(_04174_),
    .ZN(_04587_));
 AND2_X1 _29720_ (.A1(_02595_),
    .A2(_02479_),
    .ZN(_04588_));
 AND2_X1 _29721_ (.A1(_02478_),
    .A2(_02871_),
    .ZN(_04589_));
 NOR4_X1 _29722_ (.A1(_02480_),
    .A2(_04588_),
    .A3(_03893_),
    .A4(_04589_),
    .ZN(_04590_));
 AND4_X1 _29723_ (.A1(_04582_),
    .A2(_04584_),
    .A3(_04587_),
    .A4(_04590_),
    .ZN(_04591_));
 OAI21_X1 _29724_ (.A(_02581_),
    .B1(_04434_),
    .B2(_02408_),
    .ZN(_04593_));
 AND3_X1 _29725_ (.A1(_02924_),
    .A2(_02583_),
    .A3(_02554_),
    .ZN(_04594_));
 AND4_X1 _29726_ (.A1(_02557_),
    .A2(_02583_),
    .A3(_02403_),
    .A4(_02459_),
    .ZN(_04595_));
 NOR4_X1 _29727_ (.A1(_02918_),
    .A2(_04151_),
    .A3(_04594_),
    .A4(_04595_),
    .ZN(_04596_));
 OAI21_X1 _29728_ (.A(_02575_),
    .B1(_02610_),
    .B2(_03335_),
    .ZN(_04597_));
 AND3_X1 _29729_ (.A1(_04597_),
    .A2(_02929_),
    .A3(_03877_),
    .ZN(_04598_));
 NAND3_X1 _29730_ (.A1(_02450_),
    .A2(_02437_),
    .A3(_02596_),
    .ZN(_04599_));
 OAI211_X1 _29731_ (.A(_02437_),
    .B(_02583_),
    .C1(_02578_),
    .C2(_02571_),
    .ZN(_04600_));
 NAND4_X1 _29732_ (.A1(_02596_),
    .A2(_02452_),
    .A3(_02437_),
    .A4(_02454_),
    .ZN(_04601_));
 AND4_X1 _29733_ (.A1(_04599_),
    .A2(_02606_),
    .A3(_04600_),
    .A4(_04601_),
    .ZN(_04602_));
 AND4_X1 _29734_ (.A1(_04593_),
    .A2(_04596_),
    .A3(_04598_),
    .A4(_04602_),
    .ZN(_04604_));
 OAI21_X1 _29735_ (.A(_02391_),
    .B1(_02448_),
    .B2(_02897_),
    .ZN(_04605_));
 OAI21_X1 _29736_ (.A(_02461_),
    .B1(_02483_),
    .B2(_02408_),
    .ZN(_04606_));
 OAI211_X1 _29737_ (.A(_02461_),
    .B(_02394_),
    .C1(_02428_),
    .C2(_02429_),
    .ZN(_04607_));
 AND2_X1 _29738_ (.A1(_04606_),
    .A2(_04607_),
    .ZN(_04608_));
 NAND2_X1 _29739_ (.A1(_02595_),
    .A2(_02442_),
    .ZN(_04609_));
 OAI21_X1 _29740_ (.A(_02442_),
    .B1(_02450_),
    .B2(_02571_),
    .ZN(_04610_));
 AND4_X1 _29741_ (.A1(_03329_),
    .A2(_04608_),
    .A3(_04609_),
    .A4(_04610_),
    .ZN(_04611_));
 OAI21_X1 _29742_ (.A(_02391_),
    .B1(_02408_),
    .B2(_03888_),
    .ZN(_04612_));
 NOR2_X1 _29743_ (.A1(_02602_),
    .A2(_02924_),
    .ZN(_04613_));
 NOR2_X1 _29744_ (.A1(_04613_),
    .A2(_02419_),
    .ZN(_04615_));
 AND2_X1 _29745_ (.A1(_02527_),
    .A2(_02432_),
    .ZN(_04616_));
 AND2_X1 _29746_ (.A1(_02466_),
    .A2(_02432_),
    .ZN(_04617_));
 AND4_X1 _29747_ (.A1(_02438_),
    .A2(_02472_),
    .A3(_02434_),
    .A4(_02558_),
    .ZN(_04618_));
 NOR4_X1 _29748_ (.A1(_04615_),
    .A2(_04616_),
    .A3(_04617_),
    .A4(_04618_),
    .ZN(_04619_));
 AND4_X1 _29749_ (.A1(_04605_),
    .A2(_04611_),
    .A3(_04612_),
    .A4(_04619_),
    .ZN(_04620_));
 NAND4_X1 _29750_ (.A1(_04578_),
    .A2(_04591_),
    .A3(_04604_),
    .A4(_04620_),
    .ZN(_04621_));
 NOR2_X2 _29751_ (.A1(_04621_),
    .A2(_02616_),
    .ZN(_04622_));
 XOR2_X2 _29752_ (.A(_04562_),
    .B(_04622_),
    .Z(_04623_));
 AND4_X1 _29753_ (.A1(_02178_),
    .A2(_02227_),
    .A3(_02166_),
    .A4(_02161_),
    .ZN(_04624_));
 AND2_X1 _29754_ (.A1(_02238_),
    .A2(_02294_),
    .ZN(_04626_));
 AOI211_X1 _29755_ (.A(_04624_),
    .B(_04626_),
    .C1(_02328_),
    .C2(_02238_),
    .ZN(_04627_));
 OAI21_X1 _29756_ (.A(_03052_),
    .B1(_02200_),
    .B2(_02356_),
    .ZN(_04628_));
 OAI21_X1 _29757_ (.A(_03052_),
    .B1(_02252_),
    .B2(_02379_),
    .ZN(_04629_));
 AND3_X1 _29758_ (.A1(_04627_),
    .A2(_04628_),
    .A3(_04629_),
    .ZN(_04630_));
 AND2_X1 _29759_ (.A1(_03675_),
    .A2(_04273_),
    .ZN(_04631_));
 NAND2_X1 _29760_ (.A1(_02220_),
    .A2(_02288_),
    .ZN(_04632_));
 AND4_X1 _29761_ (.A1(_03672_),
    .A2(_04631_),
    .A3(_03049_),
    .A4(_04632_),
    .ZN(_04633_));
 NAND2_X1 _29762_ (.A1(_03118_),
    .A2(_02151_),
    .ZN(_04634_));
 NAND4_X1 _29763_ (.A1(_02240_),
    .A2(_02227_),
    .A3(_02301_),
    .A4(_02150_),
    .ZN(_04635_));
 NAND4_X1 _29764_ (.A1(_02225_),
    .A2(_02227_),
    .A3(_02301_),
    .A4(_02150_),
    .ZN(_04637_));
 OAI21_X1 _29765_ (.A(_02151_),
    .B1(_02221_),
    .B2(_02223_),
    .ZN(_04638_));
 AND4_X1 _29766_ (.A1(_04634_),
    .A2(_04635_),
    .A3(_04637_),
    .A4(_04638_),
    .ZN(_04639_));
 NAND3_X1 _29767_ (.A1(_02347_),
    .A2(_02171_),
    .A3(_02227_),
    .ZN(_04640_));
 NAND2_X1 _29768_ (.A1(_03448_),
    .A2(_04640_),
    .ZN(_04641_));
 AOI211_X1 _29769_ (.A(_03066_),
    .B(_04641_),
    .C1(_02239_),
    .C2(_03064_),
    .ZN(_04642_));
 AND4_X1 _29770_ (.A1(_04630_),
    .A2(_04633_),
    .A3(_04639_),
    .A4(_04642_),
    .ZN(_04643_));
 AOI221_X1 _29771_ (.A(_04259_),
    .B1(_02221_),
    .B2(_02180_),
    .C1(_02301_),
    .C2(_04260_),
    .ZN(_04644_));
 AND2_X1 _29772_ (.A1(_02358_),
    .A2(_02337_),
    .ZN(_04645_));
 INV_X1 _29773_ (.A(_04645_),
    .ZN(_04646_));
 OAI21_X1 _29774_ (.A(_02339_),
    .B1(_03056_),
    .B2(_02368_),
    .ZN(_04648_));
 OAI21_X1 _29775_ (.A(_02339_),
    .B1(_02379_),
    .B2(_02223_),
    .ZN(_04649_));
 NAND4_X1 _29776_ (.A1(_04644_),
    .A2(_04646_),
    .A3(_04648_),
    .A4(_04649_),
    .ZN(_04650_));
 NOR2_X1 _29777_ (.A1(_02376_),
    .A2(_02280_),
    .ZN(_04651_));
 NAND3_X1 _29778_ (.A1(_02167_),
    .A2(_02179_),
    .A3(_02171_),
    .ZN(_04652_));
 AND3_X1 _29779_ (.A1(_03079_),
    .A2(_04007_),
    .A3(_04652_),
    .ZN(_04653_));
 OAI21_X1 _29780_ (.A(_02326_),
    .B1(_02363_),
    .B2(_02345_),
    .ZN(_04654_));
 NAND4_X1 _29781_ (.A1(_04653_),
    .A2(_03732_),
    .A3(_03733_),
    .A4(_04654_),
    .ZN(_04655_));
 NOR4_X1 _29782_ (.A1(_04650_),
    .A2(_04651_),
    .A3(_03504_),
    .A4(_04655_),
    .ZN(_04656_));
 AND2_X1 _29783_ (.A1(_02287_),
    .A2(_02199_),
    .ZN(_04657_));
 AOI211_X1 _29784_ (.A(_04657_),
    .B(_03100_),
    .C1(_02369_),
    .C2(_04316_),
    .ZN(_04659_));
 AND2_X1 _29785_ (.A1(_02212_),
    .A2(_02214_),
    .ZN(_04660_));
 NOR4_X1 _29786_ (.A1(_03713_),
    .A2(_04660_),
    .A3(_03092_),
    .A4(_03716_),
    .ZN(_04661_));
 OAI21_X1 _29787_ (.A(_02209_),
    .B1(_02252_),
    .B2(_02194_),
    .ZN(_04662_));
 NAND2_X1 _29788_ (.A1(_02209_),
    .A2(_02356_),
    .ZN(_04663_));
 OAI211_X1 _29789_ (.A(_02284_),
    .B(_02226_),
    .C1(_02318_),
    .C2(_02294_),
    .ZN(_04664_));
 AND4_X1 _29790_ (.A1(_02372_),
    .A2(_04662_),
    .A3(_04663_),
    .A4(_04664_),
    .ZN(_04665_));
 OAI21_X1 _29791_ (.A(_02192_),
    .B1(_02345_),
    .B2(_02164_),
    .ZN(_04666_));
 NAND2_X1 _29792_ (.A1(_02192_),
    .A2(_02254_),
    .ZN(_04667_));
 AND3_X1 _29793_ (.A1(_03112_),
    .A2(_04666_),
    .A3(_04667_),
    .ZN(_04668_));
 AND4_X1 _29794_ (.A1(_04659_),
    .A2(_04661_),
    .A3(_04665_),
    .A4(_04668_),
    .ZN(_04670_));
 OAI21_X1 _29795_ (.A(_02245_),
    .B1(_02200_),
    .B2(_04316_),
    .ZN(_04671_));
 NAND4_X1 _29796_ (.A1(_02278_),
    .A2(_02239_),
    .A3(_02260_),
    .A4(_02261_),
    .ZN(_04672_));
 NAND4_X1 _29797_ (.A1(_02260_),
    .A2(_03080_),
    .A3(_02240_),
    .A4(_02261_),
    .ZN(_04673_));
 AND3_X1 _29798_ (.A1(_04671_),
    .A2(_04672_),
    .A3(_04673_),
    .ZN(_04674_));
 NAND2_X1 _29799_ (.A1(_02356_),
    .A2(_02264_),
    .ZN(_04675_));
 AND2_X1 _29800_ (.A1(_02252_),
    .A2(_02264_),
    .ZN(_04676_));
 INV_X1 _29801_ (.A(_04676_),
    .ZN(_04677_));
 NAND2_X1 _29802_ (.A1(_02254_),
    .A2(_02264_),
    .ZN(_04678_));
 OAI21_X1 _29803_ (.A(_02264_),
    .B1(_03056_),
    .B2(_02345_),
    .ZN(_04679_));
 AND4_X1 _29804_ (.A1(_04675_),
    .A2(_04677_),
    .A3(_04678_),
    .A4(_04679_),
    .ZN(_04681_));
 AOI21_X1 _29805_ (.A(_03461_),
    .B1(_04277_),
    .B2(_02205_),
    .ZN(_04682_));
 AND2_X1 _29806_ (.A1(_02345_),
    .A2(_02274_),
    .ZN(_04683_));
 AND3_X1 _29807_ (.A1(_02274_),
    .A2(_02198_),
    .A3(_02240_),
    .ZN(_04684_));
 NOR4_X1 _29808_ (.A1(_04682_),
    .A2(_03125_),
    .A3(_04683_),
    .A4(_04684_),
    .ZN(_04685_));
 AND4_X1 _29809_ (.A1(_02269_),
    .A2(_03456_),
    .A3(_03691_),
    .A4(_04313_),
    .ZN(_04686_));
 AND4_X1 _29810_ (.A1(_04674_),
    .A2(_04681_),
    .A3(_04685_),
    .A4(_04686_),
    .ZN(_04687_));
 NAND4_X1 _29811_ (.A1(_04643_),
    .A2(_04656_),
    .A3(_04670_),
    .A4(_04687_),
    .ZN(_04688_));
 NOR2_X2 _29812_ (.A1(_04688_),
    .A2(_02282_),
    .ZN(_04689_));
 XNOR2_X1 _29813_ (.A(_04385_),
    .B(_04689_),
    .ZN(_04690_));
 XNOR2_X1 _29814_ (.A(_04623_),
    .B(_04690_),
    .ZN(_04692_));
 AND2_X1 _29815_ (.A1(_02811_),
    .A2(_03952_),
    .ZN(_04693_));
 AND2_X1 _29816_ (.A1(_03558_),
    .A2(_02754_),
    .ZN(_04694_));
 NOR4_X1 _29817_ (.A1(_04693_),
    .A2(_04694_),
    .A3(_03164_),
    .A4(_04087_),
    .ZN(_04695_));
 NAND2_X1 _29818_ (.A1(_02796_),
    .A2(_02731_),
    .ZN(_04696_));
 AOI22_X1 _29819_ (.A1(_02782_),
    .A2(_02828_),
    .B1(_02831_),
    .B2(_03182_),
    .ZN(_04697_));
 NAND4_X1 _29820_ (.A1(_04695_),
    .A2(_03595_),
    .A3(_04696_),
    .A4(_04697_),
    .ZN(_04698_));
 AND3_X1 _29821_ (.A1(_02798_),
    .A2(_02822_),
    .A3(_03934_),
    .ZN(_04699_));
 AOI22_X1 _29822_ (.A1(_03952_),
    .A2(_03541_),
    .B1(_02698_),
    .B2(_02732_),
    .ZN(_04700_));
 AOI22_X1 _29823_ (.A1(_02769_),
    .A2(_02686_),
    .B1(_02823_),
    .B2(_02654_),
    .ZN(_04701_));
 NAND4_X1 _29824_ (.A1(_04699_),
    .A2(_02783_),
    .A3(_04700_),
    .A4(_04701_),
    .ZN(_04703_));
 OAI221_X1 _29825_ (.A(_02826_),
    .B1(_03200_),
    .B2(_02817_),
    .C1(_03189_),
    .C2(_03572_),
    .ZN(_04704_));
 AOI22_X1 _29826_ (.A1(_02664_),
    .A2(_02782_),
    .B1(_02654_),
    .B2(_02754_),
    .ZN(_04705_));
 NAND2_X1 _29827_ (.A1(_03169_),
    .A2(_02680_),
    .ZN(_04706_));
 OAI211_X1 _29828_ (.A(_04705_),
    .B(_04706_),
    .C1(_02776_),
    .C2(_02691_),
    .ZN(_04707_));
 NOR4_X1 _29829_ (.A1(_04698_),
    .A2(_04703_),
    .A3(_04704_),
    .A4(_04707_),
    .ZN(_04708_));
 AND2_X1 _29830_ (.A1(_02780_),
    .A2(_02632_),
    .ZN(_04709_));
 AND2_X1 _29831_ (.A1(_02664_),
    .A2(_03203_),
    .ZN(_04710_));
 AND3_X1 _29832_ (.A1(_03156_),
    .A2(_02661_),
    .A3(_02752_),
    .ZN(_04711_));
 OR4_X1 _29833_ (.A1(_04709_),
    .A2(_04710_),
    .A3(_03605_),
    .A4(_04711_),
    .ZN(_04712_));
 NAND4_X1 _29834_ (.A1(_02758_),
    .A2(_02771_),
    .A3(_02683_),
    .A4(_04487_),
    .ZN(_04714_));
 OAI21_X1 _29835_ (.A(_02635_),
    .B1(_02724_),
    .B2(_02813_),
    .ZN(_04715_));
 OAI211_X1 _29836_ (.A(_04715_),
    .B(_02760_),
    .C1(_03571_),
    .C2(_03190_),
    .ZN(_04716_));
 OAI221_X1 _29837_ (.A(_04477_),
    .B1(_03145_),
    .B2(_03190_),
    .C1(_02719_),
    .C2(_03200_),
    .ZN(_04717_));
 NOR4_X1 _29838_ (.A1(_04712_),
    .A2(_04714_),
    .A3(_04716_),
    .A4(_04717_),
    .ZN(_04718_));
 OAI21_X1 _29839_ (.A(_03172_),
    .B1(_02682_),
    .B2(_02796_),
    .ZN(_04719_));
 AOI221_X4 _29840_ (.A(_04051_),
    .B1(_02728_),
    .B2(_02663_),
    .C1(_02671_),
    .C2(_02732_),
    .ZN(_04720_));
 AND2_X1 _29841_ (.A1(_02821_),
    .A2(_02643_),
    .ZN(_04721_));
 AND3_X1 _29842_ (.A1(_02675_),
    .A2(_03211_),
    .A3(_03234_),
    .ZN(_04722_));
 NOR2_X1 _29843_ (.A1(_04721_),
    .A2(_04722_),
    .ZN(_04723_));
 AOI21_X1 _29844_ (.A(_03143_),
    .B1(_02689_),
    .B2(_03541_),
    .ZN(_04725_));
 AND4_X1 _29845_ (.A1(_04719_),
    .A2(_04720_),
    .A3(_04723_),
    .A4(_04725_),
    .ZN(_04726_));
 OAI21_X1 _29846_ (.A(_02717_),
    .B1(_03171_),
    .B2(_03574_),
    .ZN(_04727_));
 AOI21_X1 _29847_ (.A(_02700_),
    .B1(_03151_),
    .B2(_02776_),
    .ZN(_04728_));
 NOR3_X1 _29848_ (.A1(_04728_),
    .A2(_03220_),
    .A3(_04457_),
    .ZN(_04729_));
 AOI21_X1 _29849_ (.A(_03535_),
    .B1(_03152_),
    .B2(_03207_),
    .ZN(_04730_));
 AND2_X1 _29850_ (.A1(_02709_),
    .A2(_02815_),
    .ZN(_04731_));
 AND4_X1 _29851_ (.A1(_02636_),
    .A2(_02662_),
    .A3(_02674_),
    .A4(_02678_),
    .ZN(_04732_));
 NOR4_X1 _29852_ (.A1(_04730_),
    .A2(_04731_),
    .A3(_03199_),
    .A4(_04732_),
    .ZN(_04733_));
 OAI21_X1 _29853_ (.A(_02812_),
    .B1(_02809_),
    .B2(_02745_),
    .ZN(_04734_));
 AND4_X1 _29854_ (.A1(_04727_),
    .A2(_04729_),
    .A3(_04733_),
    .A4(_04734_),
    .ZN(_04736_));
 AND4_X1 _29855_ (.A1(_04708_),
    .A2(_04718_),
    .A3(_04726_),
    .A4(_04736_),
    .ZN(_04737_));
 OAI211_X1 _29856_ (.A(_03233_),
    .B(_03235_),
    .C1(_03229_),
    .C2(_03189_),
    .ZN(_04738_));
 OAI21_X1 _29857_ (.A(_03204_),
    .B1(_03160_),
    .B2(_04092_),
    .ZN(_04739_));
 OAI21_X1 _29858_ (.A(_02723_),
    .B1(_02698_),
    .B2(_03209_),
    .ZN(_04740_));
 AOI22_X1 _29859_ (.A1(_03913_),
    .A2(_02742_),
    .B1(_03169_),
    .B2(_02665_),
    .ZN(_04741_));
 NAND3_X1 _29860_ (.A1(_04739_),
    .A2(_04740_),
    .A3(_04741_),
    .ZN(_04742_));
 AND3_X1 _29861_ (.A1(_02761_),
    .A2(_03246_),
    .A3(_02678_),
    .ZN(_04743_));
 AOI211_X1 _29862_ (.A(_04738_),
    .B(_04742_),
    .C1(_02693_),
    .C2(_04743_),
    .ZN(_04744_));
 NAND2_X2 _29863_ (.A1(_04737_),
    .A2(_04744_),
    .ZN(_04745_));
 XNOR2_X1 _29864_ (.A(_04692_),
    .B(_04745_),
    .ZN(_04747_));
 XNOR2_X1 _29865_ (.A(_04747_),
    .B(_17159_),
    .ZN(_04748_));
 MUX2_X1 _29866_ (.A(_04503_),
    .B(_04748_),
    .S(_01825_),
    .Z(_00714_));
 XOR2_X1 _29867_ (.A(_17160_),
    .B(_17031_),
    .Z(_04749_));
 NAND2_X1 _29868_ (.A1(_02192_),
    .A2(_02337_),
    .ZN(_04750_));
 OAI21_X1 _29869_ (.A(_02191_),
    .B1(_02345_),
    .B2(_02268_),
    .ZN(_04751_));
 AND4_X1 _29870_ (.A1(_04750_),
    .A2(_04751_),
    .A3(_03112_),
    .A4(_03993_),
    .ZN(_04752_));
 OAI211_X1 _29871_ (.A(_02284_),
    .B(_02226_),
    .C1(_02370_),
    .C2(_02361_),
    .ZN(_04753_));
 OAI21_X1 _29872_ (.A(_02215_),
    .B1(_02216_),
    .B2(_02333_),
    .ZN(_04754_));
 NAND4_X1 _29873_ (.A1(_04752_),
    .A2(_02346_),
    .A3(_04753_),
    .A4(_04754_),
    .ZN(_04755_));
 AND2_X1 _29874_ (.A1(_02195_),
    .A2(_02350_),
    .ZN(_04757_));
 AND2_X1 _29875_ (.A1(_03699_),
    .A2(_02351_),
    .ZN(_04758_));
 AOI211_X1 _29876_ (.A(_04757_),
    .B(_04758_),
    .C1(_02223_),
    .C2(_02351_),
    .ZN(_04759_));
 NAND2_X1 _29877_ (.A1(_03699_),
    .A2(_02326_),
    .ZN(_04760_));
 OAI21_X1 _29878_ (.A(_02325_),
    .B1(_02248_),
    .B2(_02370_),
    .ZN(_04761_));
 OAI21_X1 _29879_ (.A(_02325_),
    .B1(_02216_),
    .B2(_02204_),
    .ZN(_04762_));
 AND4_X1 _29880_ (.A1(_03078_),
    .A2(_03507_),
    .A3(_04762_),
    .A4(_04652_),
    .ZN(_04763_));
 NAND4_X1 _29881_ (.A1(_04759_),
    .A2(_04760_),
    .A3(_04761_),
    .A4(_04763_),
    .ZN(_04764_));
 AND3_X1 _29882_ (.A1(_02320_),
    .A2(_02168_),
    .A3(_02171_),
    .ZN(_04765_));
 AOI211_X1 _29883_ (.A(_04765_),
    .B(_03998_),
    .C1(_02337_),
    .C2(_02173_),
    .ZN(_04766_));
 OAI21_X1 _29884_ (.A(_02212_),
    .B1(_03062_),
    .B2(_02221_),
    .ZN(_04768_));
 OAI21_X1 _29885_ (.A(_02287_),
    .B1(_03056_),
    .B2(_02345_),
    .ZN(_04769_));
 OAI21_X1 _29886_ (.A(_02287_),
    .B1(_02379_),
    .B2(_02276_),
    .ZN(_04770_));
 NAND4_X1 _29887_ (.A1(_04766_),
    .A2(_04768_),
    .A3(_04769_),
    .A4(_04770_),
    .ZN(_04771_));
 AND4_X1 _29888_ (.A1(_02296_),
    .A2(_02305_),
    .A3(_03517_),
    .A4(_03742_),
    .ZN(_04772_));
 OAI21_X1 _29889_ (.A(_02180_),
    .B1(_02379_),
    .B2(_02309_),
    .ZN(_04773_));
 OAI211_X1 _29890_ (.A(_02180_),
    .B(_02158_),
    .C1(_02162_),
    .C2(_02240_),
    .ZN(_04774_));
 NAND3_X1 _29891_ (.A1(_04772_),
    .A2(_04773_),
    .A3(_04774_),
    .ZN(_04775_));
 OR4_X1 _29892_ (.A1(_04755_),
    .A2(_04764_),
    .A3(_04771_),
    .A4(_04775_),
    .ZN(_04776_));
 NAND3_X1 _29893_ (.A1(_02248_),
    .A2(_02171_),
    .A3(_02261_),
    .ZN(_04777_));
 OAI211_X1 _29894_ (.A(_02171_),
    .B(_02261_),
    .C1(_02167_),
    .C2(_02222_),
    .ZN(_04779_));
 AND4_X1 _29895_ (.A1(_04777_),
    .A2(_04033_),
    .A3(_02256_),
    .A4(_04779_),
    .ZN(_04780_));
 OAI21_X1 _29896_ (.A(_02264_),
    .B1(_02327_),
    .B2(_02347_),
    .ZN(_04781_));
 OAI211_X1 _29897_ (.A(_02264_),
    .B(_02275_),
    .C1(_03075_),
    .C2(_02285_),
    .ZN(_04782_));
 AND4_X1 _29898_ (.A1(_04677_),
    .A2(_04780_),
    .A3(_04781_),
    .A4(_04782_),
    .ZN(_04783_));
 AND2_X1 _29899_ (.A1(_02216_),
    .A2(_02270_),
    .ZN(_04784_));
 INV_X1 _29900_ (.A(_04784_),
    .ZN(_04785_));
 INV_X1 _29901_ (.A(_03126_),
    .ZN(_04786_));
 OAI211_X1 _29902_ (.A(_02274_),
    .B(_02162_),
    .C1(_02375_),
    .C2(_02301_),
    .ZN(_04787_));
 AND4_X1 _29903_ (.A1(_04310_),
    .A2(_04785_),
    .A3(_04786_),
    .A4(_04787_),
    .ZN(_04788_));
 OAI21_X1 _29904_ (.A(_02235_),
    .B1(_02248_),
    .B2(_02370_),
    .ZN(_04790_));
 OAI211_X1 _29905_ (.A(_02235_),
    .B(_02353_),
    .C1(_03075_),
    .C2(_02285_),
    .ZN(_04791_));
 OAI221_X1 _29906_ (.A(_02235_),
    .B1(_02271_),
    .B2(_02301_),
    .C1(_03454_),
    .C2(_02225_),
    .ZN(_04792_));
 AND4_X1 _29907_ (.A1(_04788_),
    .A2(_04790_),
    .A3(_04791_),
    .A4(_04792_),
    .ZN(_04793_));
 NAND2_X1 _29908_ (.A1(_02252_),
    .A2(_02152_),
    .ZN(_04794_));
 OAI21_X1 _29909_ (.A(_02334_),
    .B1(_04286_),
    .B2(_03062_),
    .ZN(_04795_));
 OAI21_X1 _29910_ (.A(_02334_),
    .B1(_02368_),
    .B2(_02337_),
    .ZN(_04796_));
 OAI21_X1 _29911_ (.A(_02152_),
    .B1(_03118_),
    .B2(_02246_),
    .ZN(_04797_));
 AND4_X1 _29912_ (.A1(_04794_),
    .A2(_04795_),
    .A3(_04796_),
    .A4(_04797_),
    .ZN(_04798_));
 NOR2_X1 _29913_ (.A1(_03050_),
    .A2(_04280_),
    .ZN(_04799_));
 OAI221_X1 _29914_ (.A(_02220_),
    .B1(_02375_),
    .B2(_02301_),
    .C1(_02275_),
    .C2(_02225_),
    .ZN(_04801_));
 OAI21_X1 _29915_ (.A(_02238_),
    .B1(_02189_),
    .B2(_02370_),
    .ZN(_04802_));
 AND4_X1 _29916_ (.A1(_04799_),
    .A2(_04273_),
    .A3(_04801_),
    .A4(_04802_),
    .ZN(_04803_));
 NAND4_X1 _29917_ (.A1(_04783_),
    .A2(_04793_),
    .A3(_04798_),
    .A4(_04803_),
    .ZN(_04804_));
 NOR2_X2 _29918_ (.A1(_04776_),
    .A2(_04804_),
    .ZN(_04805_));
 INV_X1 _29919_ (.A(_04805_),
    .ZN(_04806_));
 XNOR2_X1 _29920_ (.A(_04562_),
    .B(_04806_),
    .ZN(_04807_));
 OAI21_X1 _29921_ (.A(_02493_),
    .B1(_03895_),
    .B2(_02511_),
    .ZN(_04808_));
 AND4_X1 _29922_ (.A1(_02387_),
    .A2(_02401_),
    .A3(_02403_),
    .A4(_02524_),
    .ZN(_04809_));
 AND2_X1 _29923_ (.A1(_02503_),
    .A2(_02570_),
    .ZN(_04810_));
 AOI211_X1 _29924_ (.A(_04809_),
    .B(_04810_),
    .C1(_02503_),
    .C2(_03895_),
    .ZN(_04812_));
 OAI21_X1 _29925_ (.A(_02503_),
    .B1(_02466_),
    .B2(_02467_),
    .ZN(_04813_));
 OAI211_X1 _29926_ (.A(_03295_),
    .B(_02524_),
    .C1(_02476_),
    .C2(_02541_),
    .ZN(_04814_));
 AND4_X1 _29927_ (.A1(_04808_),
    .A2(_04812_),
    .A3(_04813_),
    .A4(_04814_),
    .ZN(_04815_));
 OAI21_X1 _29928_ (.A(_02574_),
    .B1(_02921_),
    .B2(_02476_),
    .ZN(_04816_));
 NAND4_X1 _29929_ (.A1(_02583_),
    .A2(_02586_),
    .A3(_02609_),
    .A4(_02392_),
    .ZN(_04817_));
 OAI21_X1 _29930_ (.A(_02574_),
    .B1(_02398_),
    .B2(_02489_),
    .ZN(_04818_));
 AND3_X1 _29931_ (.A1(_04816_),
    .A2(_04817_),
    .A3(_04818_),
    .ZN(_04819_));
 OAI21_X1 _29932_ (.A(_02581_),
    .B1(_02602_),
    .B2(_02924_),
    .ZN(_04820_));
 OAI21_X1 _29933_ (.A(_02581_),
    .B1(_02467_),
    .B2(_02455_),
    .ZN(_04821_));
 AND3_X1 _29934_ (.A1(_04819_),
    .A2(_04820_),
    .A3(_04821_),
    .ZN(_04823_));
 OAI21_X1 _29935_ (.A(_02599_),
    .B1(_02420_),
    .B2(_02522_),
    .ZN(_04824_));
 OAI211_X1 _29936_ (.A(_02436_),
    .B(_02583_),
    .C1(_02570_),
    .C2(_02495_),
    .ZN(_04825_));
 OAI211_X1 _29937_ (.A(_04824_),
    .B(_04825_),
    .C1(_02932_),
    .C2(_03894_),
    .ZN(_04826_));
 NAND2_X1 _29938_ (.A1(_02547_),
    .A2(_02593_),
    .ZN(_04827_));
 NAND3_X1 _29939_ (.A1(_04827_),
    .A2(_02608_),
    .A3(_02919_),
    .ZN(_04828_));
 NOR4_X1 _29940_ (.A1(_04152_),
    .A2(_04826_),
    .A3(_02918_),
    .A4(_04828_),
    .ZN(_04829_));
 NAND4_X1 _29941_ (.A1(_02521_),
    .A2(_04172_),
    .A3(_04586_),
    .A4(_03899_),
    .ZN(_04830_));
 AOI21_X1 _29942_ (.A(_02488_),
    .B1(_02933_),
    .B2(_03883_),
    .ZN(_04831_));
 NOR4_X1 _29943_ (.A1(_04830_),
    .A2(_02900_),
    .A3(_04589_),
    .A4(_04831_),
    .ZN(_04832_));
 NAND4_X1 _29944_ (.A1(_04815_),
    .A2(_04823_),
    .A3(_04829_),
    .A4(_04832_),
    .ZN(_04834_));
 NAND2_X1 _29945_ (.A1(_02507_),
    .A2(_02442_),
    .ZN(_04835_));
 NAND2_X1 _29946_ (.A1(_04170_),
    .A2(_02461_),
    .ZN(_04836_));
 AND4_X1 _29947_ (.A1(_03333_),
    .A2(_03849_),
    .A3(_04419_),
    .A4(_04836_),
    .ZN(_04837_));
 OAI21_X1 _29948_ (.A(_02441_),
    .B1(_02404_),
    .B2(_02571_),
    .ZN(_04838_));
 OAI211_X1 _29949_ (.A(_02927_),
    .B(_02441_),
    .C1(_02926_),
    .C2(_02434_),
    .ZN(_04839_));
 AND4_X1 _29950_ (.A1(_04835_),
    .A2(_04837_),
    .A3(_04838_),
    .A4(_04839_),
    .ZN(_04840_));
 AOI21_X1 _29951_ (.A(_02885_),
    .B1(_02425_),
    .B2(_04166_),
    .ZN(_04841_));
 OAI211_X1 _29952_ (.A(_03302_),
    .B(_02890_),
    .C1(_03308_),
    .C2(_02419_),
    .ZN(_04842_));
 AOI21_X1 _29953_ (.A(_02419_),
    .B1(_02517_),
    .B2(_02447_),
    .ZN(_04843_));
 NAND2_X1 _29954_ (.A1(_04133_),
    .A2(_04134_),
    .ZN(_04845_));
 NOR4_X1 _29955_ (.A1(_04841_),
    .A2(_04842_),
    .A3(_04843_),
    .A4(_04845_),
    .ZN(_04846_));
 NAND2_X1 _29956_ (.A1(_02560_),
    .A2(_02466_),
    .ZN(_04847_));
 AND3_X1 _29957_ (.A1(_02533_),
    .A2(_02926_),
    .A3(_02927_),
    .ZN(_04848_));
 AOI21_X1 _29958_ (.A(_04848_),
    .B1(_02534_),
    .B2(_02921_),
    .ZN(_04849_));
 OAI21_X1 _29959_ (.A(_02560_),
    .B1(_02448_),
    .B2(_02398_),
    .ZN(_04850_));
 OAI21_X1 _29960_ (.A(_02533_),
    .B1(_02500_),
    .B2(_02871_),
    .ZN(_04851_));
 AND4_X1 _29961_ (.A1(_04847_),
    .A2(_04849_),
    .A3(_04850_),
    .A4(_04851_),
    .ZN(_04852_));
 NAND2_X1 _29962_ (.A1(_02540_),
    .A2(_02466_),
    .ZN(_04853_));
 OAI21_X1 _29963_ (.A(_02540_),
    .B1(_02410_),
    .B2(_02481_),
    .ZN(_04854_));
 NAND4_X1 _29964_ (.A1(_03321_),
    .A2(_04853_),
    .A3(_04576_),
    .A4(_04854_),
    .ZN(_04856_));
 NOR4_X1 _29965_ (.A1(_04856_),
    .A2(_04394_),
    .A3(_02550_),
    .A4(_04564_),
    .ZN(_04857_));
 NAND4_X1 _29966_ (.A1(_04840_),
    .A2(_04846_),
    .A3(_04852_),
    .A4(_04857_),
    .ZN(_04858_));
 NOR2_X1 _29967_ (.A1(_04834_),
    .A2(_04858_),
    .ZN(_04859_));
 INV_X2 _29968_ (.A(_04859_),
    .ZN(_04860_));
 XNOR2_X2 _29969_ (.A(_02139_),
    .B(_04860_),
    .ZN(_04861_));
 XNOR2_X1 _29970_ (.A(_04807_),
    .B(_04861_),
    .ZN(_04862_));
 AND2_X1 _29971_ (.A1(_02828_),
    .A2(_02813_),
    .ZN(_04863_));
 NAND2_X1 _29972_ (.A1(_04074_),
    .A2(_02822_),
    .ZN(_04864_));
 OR4_X1 _29973_ (.A1(_04863_),
    .A2(_04864_),
    .A3(_04721_),
    .A4(_03594_),
    .ZN(_04865_));
 AND3_X1 _29974_ (.A1(_02675_),
    .A2(_02676_),
    .A3(_03211_),
    .ZN(_04867_));
 AND2_X1 _29975_ (.A1(_02811_),
    .A2(_02704_),
    .ZN(_04868_));
 AOI211_X1 _29976_ (.A(_04867_),
    .B(_04868_),
    .C1(_02811_),
    .C2(_04092_),
    .ZN(_04869_));
 OAI221_X1 _29977_ (.A(_04869_),
    .B1(_02638_),
    .B2(_03914_),
    .C1(_03603_),
    .C2(_04468_),
    .ZN(_04870_));
 AOI21_X1 _29978_ (.A(_03200_),
    .B1(_03157_),
    .B2(_02817_),
    .ZN(_04871_));
 OR4_X1 _29979_ (.A1(_03916_),
    .A2(_04871_),
    .A3(_03608_),
    .A4(_04451_),
    .ZN(_04872_));
 AOI21_X1 _29980_ (.A(_03189_),
    .B1(_03145_),
    .B2(_02816_),
    .ZN(_04873_));
 OAI21_X1 _29981_ (.A(_02826_),
    .B1(_03189_),
    .B2(_03207_),
    .ZN(_04874_));
 AND4_X1 _29982_ (.A1(_02761_),
    .A2(_02823_),
    .A3(_02743_),
    .A4(_02656_),
    .ZN(_04875_));
 OR4_X1 _29983_ (.A1(_04722_),
    .A2(_04873_),
    .A3(_04874_),
    .A4(_04875_),
    .ZN(_04876_));
 NOR4_X1 _29984_ (.A1(_04865_),
    .A2(_04870_),
    .A3(_04872_),
    .A4(_04876_),
    .ZN(_04878_));
 AND2_X1 _29985_ (.A1(_02732_),
    .A2(_02647_),
    .ZN(_04879_));
 OAI211_X1 _29986_ (.A(_03181_),
    .B(_04109_),
    .C1(_03152_),
    .C2(_03535_),
    .ZN(_04880_));
 NAND2_X1 _29987_ (.A1(_02724_),
    .A2(_02742_),
    .ZN(_04881_));
 NAND2_X1 _29988_ (.A1(_02738_),
    .A2(_04881_),
    .ZN(_04882_));
 OAI211_X1 _29989_ (.A(_04696_),
    .B(_04106_),
    .C1(_04496_),
    .C2(_02829_),
    .ZN(_04883_));
 OR4_X1 _29990_ (.A1(_04879_),
    .A2(_04880_),
    .A3(_04882_),
    .A4(_04883_),
    .ZN(_04884_));
 AND2_X1 _29991_ (.A1(_03175_),
    .A2(_03197_),
    .ZN(_04885_));
 AND2_X1 _29992_ (.A1(_02695_),
    .A2(_02658_),
    .ZN(_04886_));
 NAND2_X1 _29993_ (.A1(_02670_),
    .A2(_02695_),
    .ZN(_04887_));
 NAND3_X1 _29994_ (.A1(_04887_),
    .A2(_03543_),
    .A3(_02705_),
    .ZN(_04889_));
 AOI21_X1 _29995_ (.A(_02700_),
    .B1(_02715_),
    .B2(_02688_),
    .ZN(_04890_));
 NOR2_X1 _29996_ (.A1(_02700_),
    .A2(_03229_),
    .ZN(_04891_));
 OR4_X1 _29997_ (.A1(_04886_),
    .A2(_04889_),
    .A3(_04890_),
    .A4(_04891_),
    .ZN(_04892_));
 NOR4_X1 _29998_ (.A1(_04884_),
    .A2(_04885_),
    .A3(_03973_),
    .A4(_04892_),
    .ZN(_04893_));
 INV_X1 _29999_ (.A(_02631_),
    .ZN(_04894_));
 NAND2_X1 _30000_ (.A1(_02635_),
    .A2(_03237_),
    .ZN(_04895_));
 NAND4_X1 _30001_ (.A1(_04894_),
    .A2(_02655_),
    .A3(_02644_),
    .A4(_04895_),
    .ZN(_04896_));
 INV_X1 _30002_ (.A(_03586_),
    .ZN(_04897_));
 NAND2_X1 _30003_ (.A1(_02717_),
    .A2(_03209_),
    .ZN(_04898_));
 NAND4_X1 _30004_ (.A1(_04897_),
    .A2(_04898_),
    .A3(_03248_),
    .A4(_04099_),
    .ZN(_04900_));
 OAI211_X1 _30005_ (.A(_02662_),
    .B(_02622_),
    .C1(_03952_),
    .C2(_02696_),
    .ZN(_04901_));
 NAND2_X1 _30006_ (.A1(_02665_),
    .A2(_02658_),
    .ZN(_04902_));
 NAND2_X1 _30007_ (.A1(_02664_),
    .A2(_02765_),
    .ZN(_04903_));
 NAND4_X1 _30008_ (.A1(_03249_),
    .A2(_04901_),
    .A3(_04902_),
    .A4(_04903_),
    .ZN(_04904_));
 OAI21_X1 _30009_ (.A(_02723_),
    .B1(_02641_),
    .B2(_04092_),
    .ZN(_04905_));
 OAI21_X1 _30010_ (.A(_04905_),
    .B1(_03155_),
    .B2(_03146_),
    .ZN(_04906_));
 NOR4_X1 _30011_ (.A1(_04896_),
    .A2(_04900_),
    .A3(_04904_),
    .A4(_04906_),
    .ZN(_04907_));
 NAND2_X1 _30012_ (.A1(_02796_),
    .A2(_03172_),
    .ZN(_04908_));
 NAND4_X1 _30013_ (.A1(_03908_),
    .A2(_02771_),
    .A3(_04060_),
    .A4(_04908_),
    .ZN(_04909_));
 NAND2_X1 _30014_ (.A1(_03558_),
    .A2(_03204_),
    .ZN(_04911_));
 OAI21_X1 _30015_ (.A(_03204_),
    .B1(_02654_),
    .B2(_02724_),
    .ZN(_04912_));
 NAND4_X1 _30016_ (.A1(_02787_),
    .A2(_03554_),
    .A3(_04911_),
    .A4(_04912_),
    .ZN(_04913_));
 OAI21_X1 _30017_ (.A(_02799_),
    .B1(_02641_),
    .B2(_04092_),
    .ZN(_04914_));
 OAI21_X1 _30018_ (.A(_02799_),
    .B1(_03952_),
    .B2(_02793_),
    .ZN(_04915_));
 NAND4_X1 _30019_ (.A1(_02694_),
    .A2(_02748_),
    .A3(_02829_),
    .A4(_02752_),
    .ZN(_04916_));
 NAND3_X1 _30020_ (.A1(_04914_),
    .A2(_04915_),
    .A3(_04916_),
    .ZN(_04917_));
 OAI21_X1 _30021_ (.A(_02759_),
    .B1(_02641_),
    .B2(_03182_),
    .ZN(_04918_));
 OAI211_X1 _30022_ (.A(_02754_),
    .B(_02748_),
    .C1(_02652_),
    .C2(_03528_),
    .ZN(_04919_));
 NAND3_X1 _30023_ (.A1(_04918_),
    .A2(_03567_),
    .A3(_04919_),
    .ZN(_04920_));
 NOR4_X1 _30024_ (.A1(_04909_),
    .A2(_04913_),
    .A3(_04917_),
    .A4(_04920_),
    .ZN(_04922_));
 NAND4_X1 _30025_ (.A1(_04878_),
    .A2(_04893_),
    .A3(_04907_),
    .A4(_04922_),
    .ZN(_04923_));
 NOR2_X2 _30026_ (.A1(_04923_),
    .A2(_03199_),
    .ZN(_04924_));
 XNOR2_X1 _30027_ (.A(_04862_),
    .B(_04924_),
    .ZN(_04925_));
 XNOR2_X1 _30028_ (.A(_04925_),
    .B(_17160_),
    .ZN(_04926_));
 MUX2_X1 _30029_ (.A(_04749_),
    .B(_04926_),
    .S(_01825_),
    .Z(_00715_));
 XOR2_X1 _30030_ (.A(_17161_),
    .B(_17032_),
    .Z(_04927_));
 XNOR2_X1 _30031_ (.A(_04805_),
    .B(_01037_),
    .ZN(_04928_));
 XOR2_X1 _30032_ (.A(_04928_),
    .B(_03253_),
    .Z(_04929_));
 XNOR2_X1 _30033_ (.A(_02050_),
    .B(_02617_),
    .ZN(_04930_));
 XNOR2_X1 _30034_ (.A(_04929_),
    .B(_04930_),
    .ZN(_04932_));
 BUF_X2 _30035_ (.A(_09038_),
    .Z(_04933_));
 MUX2_X1 _30036_ (.A(_04927_),
    .B(_04932_),
    .S(_04933_),
    .Z(_00676_));
 XOR2_X1 _30037_ (.A(_17162_),
    .B(_17033_),
    .Z(_04934_));
 XNOR2_X2 _30038_ (.A(_04806_),
    .B(_02385_),
    .ZN(_04935_));
 XNOR2_X1 _30039_ (.A(_04935_),
    .B(_03615_),
    .ZN(_04936_));
 XNOR2_X1 _30040_ (.A(_03253_),
    .B(_03043_),
    .ZN(_04937_));
 XNOR2_X1 _30041_ (.A(_04936_),
    .B(_04937_),
    .ZN(_04938_));
 XOR2_X1 _30042_ (.A(_04938_),
    .B(_17162_),
    .Z(_04939_));
 MUX2_X1 _30043_ (.A(_04934_),
    .B(_04939_),
    .S(_04933_),
    .Z(_00677_));
 XOR2_X1 _30044_ (.A(_17132_),
    .B(_17034_),
    .Z(_04941_));
 XNOR2_X1 _30045_ (.A(_03447_),
    .B(_03982_),
    .ZN(_04942_));
 XOR2_X2 _30046_ (.A(_03139_),
    .B(_03615_),
    .Z(_04943_));
 XNOR2_X1 _30047_ (.A(_04942_),
    .B(_04943_),
    .ZN(_04944_));
 XOR2_X1 _30048_ (.A(_04944_),
    .B(_17132_),
    .Z(_04945_));
 MUX2_X1 _30049_ (.A(_04941_),
    .B(_04945_),
    .S(_04933_),
    .Z(_00678_));
 XOR2_X1 _30050_ (.A(_17133_),
    .B(_17035_),
    .Z(_04946_));
 XNOR2_X1 _30051_ (.A(_04805_),
    .B(_03524_),
    .ZN(_04947_));
 XNOR2_X1 _30052_ (.A(_04947_),
    .B(_04112_),
    .ZN(_04948_));
 XNOR2_X1 _30053_ (.A(_04948_),
    .B(_03984_),
    .ZN(_04949_));
 XNOR2_X1 _30054_ (.A(_04949_),
    .B(_17133_),
    .ZN(_04951_));
 MUX2_X1 _30055_ (.A(_04946_),
    .B(_04951_),
    .S(_04933_),
    .Z(_00679_));
 XOR2_X1 _30056_ (.A(_17134_),
    .B(_17036_),
    .Z(_04952_));
 XNOR2_X2 _30057_ (.A(_04805_),
    .B(_03746_),
    .ZN(_04953_));
 XOR2_X1 _30058_ (.A(_04953_),
    .B(_04500_),
    .Z(_04954_));
 XNOR2_X1 _30059_ (.A(_04954_),
    .B(_04250_),
    .ZN(_04955_));
 XOR2_X1 _30060_ (.A(_04955_),
    .B(_17134_),
    .Z(_04956_));
 MUX2_X1 _30061_ (.A(_04952_),
    .B(_04956_),
    .S(_04933_),
    .Z(_00680_));
 XOR2_X1 _30062_ (.A(_17135_),
    .B(_17037_),
    .Z(_04957_));
 XNOR2_X1 _30063_ (.A(_04500_),
    .B(_04046_),
    .ZN(_04958_));
 XNOR2_X1 _30064_ (.A(_04446_),
    .B(_04958_),
    .ZN(_04960_));
 XNOR2_X1 _30065_ (.A(_04960_),
    .B(_04745_),
    .ZN(_04961_));
 INV_X1 _30066_ (.A(_17135_),
    .ZN(_04962_));
 XNOR2_X1 _30067_ (.A(_04961_),
    .B(_04962_),
    .ZN(_04963_));
 MUX2_X1 _30068_ (.A(_04957_),
    .B(_04963_),
    .S(_04933_),
    .Z(_00681_));
 XOR2_X1 _30069_ (.A(_17136_),
    .B(_17038_),
    .Z(_04964_));
 XOR2_X2 _30070_ (.A(_04323_),
    .B(_04745_),
    .Z(_04965_));
 XNOR2_X1 _30071_ (.A(_04623_),
    .B(_04965_),
    .ZN(_04966_));
 XNOR2_X1 _30072_ (.A(_04966_),
    .B(_04924_),
    .ZN(_04967_));
 XNOR2_X1 _30073_ (.A(_04967_),
    .B(_17136_),
    .ZN(_04968_));
 MUX2_X1 _30074_ (.A(_04964_),
    .B(_04968_),
    .S(_04933_),
    .Z(_00682_));
 XOR2_X1 _30075_ (.A(_17137_),
    .B(_17039_),
    .Z(_04970_));
 XOR2_X2 _30076_ (.A(_04924_),
    .B(_04689_),
    .Z(_04971_));
 XNOR2_X1 _30077_ (.A(_04971_),
    .B(_04861_),
    .ZN(_04972_));
 XNOR2_X1 _30078_ (.A(_04972_),
    .B(_02837_),
    .ZN(_04973_));
 XOR2_X1 _30079_ (.A(_04973_),
    .B(_17137_),
    .Z(_04974_));
 MUX2_X1 _30080_ (.A(_04970_),
    .B(_04974_),
    .S(_04933_),
    .Z(_00683_));
 XOR2_X1 _30081_ (.A(_17138_),
    .B(_17041_),
    .Z(_04975_));
 XNOR2_X1 _30082_ (.A(_04935_),
    .B(_01038_),
    .ZN(_04976_));
 XNOR2_X1 _30083_ (.A(_02050_),
    .B(_03252_),
    .ZN(_04977_));
 XNOR2_X1 _30084_ (.A(_04977_),
    .B(_04860_),
    .ZN(_04979_));
 XNOR2_X1 _30085_ (.A(_04976_),
    .B(_04979_),
    .ZN(_04980_));
 MUX2_X1 _30086_ (.A(_04975_),
    .B(_04980_),
    .S(_04933_),
    .Z(_00644_));
 XOR2_X1 _30087_ (.A(_17139_),
    .B(_17042_),
    .Z(_04981_));
 XNOR2_X1 _30088_ (.A(_04935_),
    .B(_04943_),
    .ZN(_04982_));
 XNOR2_X1 _30089_ (.A(_02617_),
    .B(_04860_),
    .ZN(_04983_));
 INV_X1 _30090_ (.A(_01039_),
    .ZN(_04984_));
 XNOR2_X1 _30091_ (.A(_03042_),
    .B(_04984_),
    .ZN(_04985_));
 XOR2_X1 _30092_ (.A(_04983_),
    .B(_04985_),
    .Z(_04986_));
 XNOR2_X1 _30093_ (.A(_04982_),
    .B(_04986_),
    .ZN(_04987_));
 MUX2_X1 _30094_ (.A(_04981_),
    .B(_04987_),
    .S(_04933_),
    .Z(_00645_));
 XOR2_X1 _30095_ (.A(_03446_),
    .B(_03524_),
    .Z(_04989_));
 XNOR2_X1 _30096_ (.A(_04989_),
    .B(_03982_),
    .ZN(_04990_));
 XNOR2_X1 _30097_ (.A(_03139_),
    .B(_02963_),
    .ZN(_04991_));
 OAI21_X1 _30098_ (.A(_09038_),
    .B1(_04990_),
    .B2(_04991_),
    .ZN(_04992_));
 AOI21_X1 _30099_ (.A(_04992_),
    .B1(_04990_),
    .B2(_04991_),
    .ZN(_04993_));
 AND2_X1 _30100_ (.A1(_01331_),
    .A2(_17043_),
    .ZN(_04994_));
 NOR2_X1 _30101_ (.A1(_04993_),
    .A2(_04994_),
    .ZN(_04995_));
 XNOR2_X1 _30102_ (.A(_04995_),
    .B(_17140_),
    .ZN(_00646_));
 XOR2_X1 _30103_ (.A(_17141_),
    .B(_17044_),
    .Z(_04996_));
 XNOR2_X1 _30104_ (.A(_04112_),
    .B(_03524_),
    .ZN(_04998_));
 XNOR2_X1 _30105_ (.A(_04953_),
    .B(_04998_),
    .ZN(_04999_));
 XNOR2_X1 _30106_ (.A(_03372_),
    .B(_04859_),
    .ZN(_05000_));
 XNOR2_X1 _30107_ (.A(_05000_),
    .B(_03821_),
    .ZN(_05001_));
 XNOR2_X1 _30108_ (.A(_04999_),
    .B(_05001_),
    .ZN(_05002_));
 XNOR2_X1 _30109_ (.A(_05002_),
    .B(_17141_),
    .ZN(_05003_));
 BUF_X2 _30110_ (.A(_09038_),
    .Z(_05004_));
 MUX2_X1 _30111_ (.A(_04996_),
    .B(_05003_),
    .S(_05004_),
    .Z(_00647_));
 XOR2_X1 _30112_ (.A(_17143_),
    .B(_17045_),
    .Z(_05005_));
 XNOR2_X1 _30113_ (.A(_04953_),
    .B(_04046_),
    .ZN(_05006_));
 XNOR2_X1 _30114_ (.A(_03902_),
    .B(_04860_),
    .ZN(_05008_));
 XNOR2_X1 _30115_ (.A(_05008_),
    .B(_04248_),
    .ZN(_05009_));
 XNOR2_X1 _30116_ (.A(_05006_),
    .B(_05009_),
    .ZN(_05010_));
 XNOR2_X1 _30117_ (.A(_05010_),
    .B(_04500_),
    .ZN(_05011_));
 XOR2_X1 _30118_ (.A(_05011_),
    .B(_17143_),
    .Z(_05012_));
 MUX2_X1 _30119_ (.A(_05005_),
    .B(_05012_),
    .S(_05004_),
    .Z(_00648_));
 XOR2_X1 _30120_ (.A(_17144_),
    .B(_17046_),
    .Z(_05013_));
 INV_X1 _30121_ (.A(_01040_),
    .ZN(_05014_));
 XNOR2_X1 _30122_ (.A(_04385_),
    .B(_05014_),
    .ZN(_05015_));
 XOR2_X1 _30123_ (.A(_05015_),
    .B(_04046_),
    .Z(_05016_));
 XNOR2_X1 _30124_ (.A(_04965_),
    .B(_04184_),
    .ZN(_05018_));
 XNOR2_X1 _30125_ (.A(_05016_),
    .B(_05018_),
    .ZN(_05019_));
 MUX2_X1 _30126_ (.A(_05013_),
    .B(_05019_),
    .S(_05004_),
    .Z(_00649_));
 XOR2_X1 _30127_ (.A(_17145_),
    .B(_17047_),
    .Z(_05020_));
 XNOR2_X1 _30128_ (.A(_04323_),
    .B(_01041_),
    .ZN(_05021_));
 XOR2_X1 _30129_ (.A(_05021_),
    .B(_04562_),
    .Z(_05022_));
 XNOR2_X1 _30130_ (.A(_04971_),
    .B(_04445_),
    .ZN(_05023_));
 XNOR2_X1 _30131_ (.A(_05022_),
    .B(_05023_),
    .ZN(_05024_));
 MUX2_X1 _30132_ (.A(_05020_),
    .B(_05024_),
    .S(_05004_),
    .Z(_00650_));
 XOR2_X1 _30133_ (.A(_17146_),
    .B(_17048_),
    .Z(_05025_));
 XOR2_X1 _30134_ (.A(_04622_),
    .B(_02139_),
    .Z(_05027_));
 XNOR2_X1 _30135_ (.A(_04805_),
    .B(_04689_),
    .ZN(_05028_));
 XNOR2_X1 _30136_ (.A(_05027_),
    .B(_05028_),
    .ZN(_05029_));
 XNOR2_X1 _30137_ (.A(_05029_),
    .B(_02837_),
    .ZN(_05030_));
 XNOR2_X1 _30138_ (.A(_05030_),
    .B(_17146_),
    .ZN(_05031_));
 MUX2_X1 _30139_ (.A(_05025_),
    .B(_05031_),
    .S(_05004_),
    .Z(_00651_));
 XOR2_X1 _30140_ (.A(_17147_),
    .B(_17049_),
    .Z(_05032_));
 XNOR2_X1 _30141_ (.A(_02617_),
    .B(_01042_),
    .ZN(_05033_));
 XNOR2_X1 _30142_ (.A(_05033_),
    .B(_04861_),
    .ZN(_05034_));
 XNOR2_X1 _30143_ (.A(_02385_),
    .B(_03252_),
    .ZN(_05035_));
 XNOR2_X1 _30144_ (.A(_05034_),
    .B(_05035_),
    .ZN(_05037_));
 MUX2_X1 _30145_ (.A(_05032_),
    .B(_05037_),
    .S(_05004_),
    .Z(_00612_));
 XOR2_X1 _30146_ (.A(_17148_),
    .B(_17050_),
    .Z(_05038_));
 XOR2_X1 _30147_ (.A(_02140_),
    .B(_04983_),
    .Z(_05039_));
 XNOR2_X1 _30148_ (.A(_04991_),
    .B(_03615_),
    .ZN(_05040_));
 XNOR2_X1 _30149_ (.A(_05039_),
    .B(_05040_),
    .ZN(_05041_));
 INV_X1 _30150_ (.A(_01043_),
    .ZN(_05042_));
 XNOR2_X1 _30151_ (.A(_05041_),
    .B(_05042_),
    .ZN(_05043_));
 MUX2_X1 _30152_ (.A(_05038_),
    .B(_05043_),
    .S(_05004_),
    .Z(_00613_));
 XOR2_X1 _30153_ (.A(_17149_),
    .B(_17052_),
    .Z(_05044_));
 XNOR2_X1 _30154_ (.A(_03372_),
    .B(_03524_),
    .ZN(_05046_));
 XNOR2_X1 _30155_ (.A(_03043_),
    .B(_05046_),
    .ZN(_05047_));
 XNOR2_X1 _30156_ (.A(_05047_),
    .B(_03982_),
    .ZN(_05048_));
 XNOR2_X1 _30157_ (.A(_05048_),
    .B(_01658_),
    .ZN(_05049_));
 MUX2_X1 _30158_ (.A(_05044_),
    .B(_05049_),
    .S(_05004_),
    .Z(_00614_));
 XOR2_X1 _30159_ (.A(_17150_),
    .B(_17053_),
    .Z(_05050_));
 XOR2_X1 _30160_ (.A(_04112_),
    .B(_03902_),
    .Z(_05051_));
 XNOR2_X1 _30161_ (.A(_03670_),
    .B(_05051_),
    .ZN(_05052_));
 XNOR2_X1 _30162_ (.A(_05000_),
    .B(_03746_),
    .ZN(_05053_));
 XNOR2_X1 _30163_ (.A(_05052_),
    .B(_05053_),
    .ZN(_05054_));
 XNOR2_X1 _30164_ (.A(_05054_),
    .B(_17150_),
    .ZN(_05056_));
 MUX2_X1 _30165_ (.A(_05050_),
    .B(_05056_),
    .S(_05004_),
    .Z(_00615_));
 XOR2_X1 _30166_ (.A(_17151_),
    .B(_17054_),
    .Z(_05057_));
 XNOR2_X1 _30167_ (.A(_03988_),
    .B(_05008_),
    .ZN(_05058_));
 XNOR2_X1 _30168_ (.A(_04184_),
    .B(_04046_),
    .ZN(_05059_));
 XNOR2_X1 _30169_ (.A(_05059_),
    .B(_04500_),
    .ZN(_05060_));
 XNOR2_X1 _30170_ (.A(_05058_),
    .B(_05060_),
    .ZN(_05061_));
 XNOR2_X1 _30171_ (.A(_05061_),
    .B(_17151_),
    .ZN(_05062_));
 MUX2_X1 _30172_ (.A(_05057_),
    .B(_05062_),
    .S(_05004_),
    .Z(_00616_));
 XOR2_X1 _30173_ (.A(_17152_),
    .B(_17055_),
    .Z(_05063_));
 XOR2_X1 _30174_ (.A(_04445_),
    .B(_01044_),
    .Z(_05065_));
 XNOR2_X1 _30175_ (.A(_05065_),
    .B(_04323_),
    .ZN(_05066_));
 XNOR2_X1 _30176_ (.A(_04249_),
    .B(_04745_),
    .ZN(_05067_));
 XNOR2_X1 _30177_ (.A(_05066_),
    .B(_05067_),
    .ZN(_05068_));
 BUF_X2 _30178_ (.A(_09038_),
    .Z(_05069_));
 MUX2_X1 _30179_ (.A(_05063_),
    .B(_05068_),
    .S(_05069_),
    .Z(_00617_));
 INV_X1 _30180_ (.A(_16678_),
    .ZN(_05070_));
 NOR2_X1 _30181_ (.A1(_01200_),
    .A2(_01201_),
    .ZN(_05071_));
 NOR2_X1 _30182_ (.A1(_01330_),
    .A2(_01199_),
    .ZN(_05072_));
 AOI221_X4 _30183_ (.A(_05070_),
    .B1(_03933_),
    .B2(_01198_),
    .C1(_05071_),
    .C2(_05072_),
    .ZN(_00599_));
 NOR3_X1 _30184_ (.A1(_01198_),
    .A2(_01199_),
    .A3(_01045_),
    .ZN(_05074_));
 INV_X1 _30185_ (.A(_05071_),
    .ZN(_05075_));
 NOR2_X1 _30186_ (.A1(_01198_),
    .A2(_01199_),
    .ZN(_05076_));
 AOI21_X1 _30187_ (.A(_05074_),
    .B1(_05075_),
    .B2(_05076_),
    .ZN(_05077_));
 AOI21_X1 _30188_ (.A(_03847_),
    .B1(_01198_),
    .B2(_01199_),
    .ZN(_05078_));
 AOI21_X1 _30189_ (.A(_05070_),
    .B1(_05077_),
    .B2(_05078_),
    .ZN(_00600_));
 AND2_X1 _30190_ (.A1(_05075_),
    .A2(_05076_),
    .ZN(_05079_));
 INV_X1 _30191_ (.A(_01046_),
    .ZN(_05080_));
 OAI211_X1 _30192_ (.A(_03749_),
    .B(_16678_),
    .C1(_05079_),
    .C2(_05080_),
    .ZN(_05081_));
 AOI21_X1 _30193_ (.A(_05081_),
    .B1(_05080_),
    .B2(_05079_),
    .ZN(_00601_));
 INV_X1 _30194_ (.A(_01200_),
    .ZN(_05083_));
 NAND3_X1 _30195_ (.A1(_05076_),
    .A2(_05083_),
    .A3(_01201_),
    .ZN(_05084_));
 INV_X1 _30196_ (.A(_01047_),
    .ZN(_05085_));
 OR2_X1 _30197_ (.A1(_05084_),
    .A2(_05085_),
    .ZN(_05086_));
 AOI21_X1 _30198_ (.A(_03847_),
    .B1(_05084_),
    .B2(_05085_),
    .ZN(_05087_));
 AOI21_X1 _30199_ (.A(_05070_),
    .B1(_05086_),
    .B2(_05087_),
    .ZN(_00602_));
 XOR2_X1 _30200_ (.A(_17154_),
    .B(_17056_),
    .Z(_05088_));
 XNOR2_X1 _30201_ (.A(_04924_),
    .B(_01048_),
    .ZN(_05089_));
 XNOR2_X1 _30202_ (.A(_04446_),
    .B(_05089_),
    .ZN(_05090_));
 XOR2_X1 _30203_ (.A(_04689_),
    .B(_04622_),
    .Z(_05091_));
 XNOR2_X1 _30204_ (.A(_05090_),
    .B(_05091_),
    .ZN(_05093_));
 MUX2_X1 _30205_ (.A(_05088_),
    .B(_05093_),
    .S(_05069_),
    .Z(_00618_));
 MUX2_X1 _30206_ (.A(_16935_),
    .B(_16807_),
    .S(_03847_),
    .Z(_00732_));
 BUF_X2 _30207_ (.A(_03836_),
    .Z(_05094_));
 MUX2_X1 _30208_ (.A(_16974_),
    .B(_16846_),
    .S(_05094_),
    .Z(_00771_));
 MUX2_X1 _30209_ (.A(_16985_),
    .B(_16857_),
    .S(_05094_),
    .Z(_00782_));
 MUX2_X1 _30210_ (.A(_16996_),
    .B(_16868_),
    .S(_05094_),
    .Z(_00793_));
 MUX2_X1 _30211_ (.A(_17007_),
    .B(_16879_),
    .S(_05094_),
    .Z(_00804_));
 MUX2_X1 _30212_ (.A(_17018_),
    .B(_16890_),
    .S(_05094_),
    .Z(_00815_));
 XOR2_X1 _30213_ (.A(_17155_),
    .B(_17057_),
    .Z(_05095_));
 XNOR2_X1 _30214_ (.A(_04805_),
    .B(_04860_),
    .ZN(_05097_));
 XNOR2_X1 _30215_ (.A(_05097_),
    .B(_02837_),
    .ZN(_05098_));
 XOR2_X1 _30216_ (.A(_05098_),
    .B(_04623_),
    .Z(_05099_));
 XNOR2_X1 _30217_ (.A(_05099_),
    .B(_17155_),
    .ZN(_05100_));
 MUX2_X1 _30218_ (.A(_05095_),
    .B(_05100_),
    .S(_05069_),
    .Z(_00619_));
 MUX2_X1 _30219_ (.A(_17029_),
    .B(_16901_),
    .S(_05094_),
    .Z(_00826_));
 MUX2_X1 _30220_ (.A(_17040_),
    .B(_16912_),
    .S(_05094_),
    .Z(_00837_));
 MUX2_X1 _30221_ (.A(_17051_),
    .B(_16923_),
    .S(_05094_),
    .Z(_00848_));
 MUX2_X1 _30222_ (.A(_17062_),
    .B(_16934_),
    .S(_05094_),
    .Z(_00859_));
 MUX2_X1 _30223_ (.A(_16946_),
    .B(_16818_),
    .S(_05094_),
    .Z(_00743_));
 BUF_X2 _30224_ (.A(_03836_),
    .Z(_05102_));
 MUX2_X1 _30225_ (.A(_16957_),
    .B(_16829_),
    .S(_05102_),
    .Z(_00754_));
 MUX2_X1 _30226_ (.A(_16966_),
    .B(_16838_),
    .S(_05102_),
    .Z(_00763_));
 MUX2_X1 _30227_ (.A(_16967_),
    .B(_16839_),
    .S(_05102_),
    .Z(_00764_));
 MUX2_X1 _30228_ (.A(_16968_),
    .B(_16840_),
    .S(_05102_),
    .Z(_00765_));
 MUX2_X1 _30229_ (.A(_16969_),
    .B(_16841_),
    .S(_05102_),
    .Z(_00766_));
 MUX2_X1 _30230_ (.A(_16970_),
    .B(_16842_),
    .S(_05102_),
    .Z(_00767_));
 MUX2_X1 _30231_ (.A(_16971_),
    .B(_16843_),
    .S(_05102_),
    .Z(_00768_));
 MUX2_X1 _30232_ (.A(_16972_),
    .B(_16844_),
    .S(_05102_),
    .Z(_00769_));
 MUX2_X1 _30233_ (.A(_16973_),
    .B(_16845_),
    .S(_05102_),
    .Z(_00770_));
 MUX2_X1 _30234_ (.A(_16975_),
    .B(_16847_),
    .S(_05102_),
    .Z(_00772_));
 BUF_X2 _30235_ (.A(_01330_),
    .Z(_05104_));
 BUF_X2 _30236_ (.A(_05104_),
    .Z(_05105_));
 MUX2_X1 _30237_ (.A(_16976_),
    .B(_16848_),
    .S(_05105_),
    .Z(_00773_));
 MUX2_X1 _30238_ (.A(_16977_),
    .B(_16849_),
    .S(_05105_),
    .Z(_00774_));
 MUX2_X1 _30239_ (.A(_16978_),
    .B(_16850_),
    .S(_05105_),
    .Z(_00775_));
 MUX2_X1 _30240_ (.A(_16979_),
    .B(_16851_),
    .S(_05105_),
    .Z(_00776_));
 MUX2_X1 _30241_ (.A(_16980_),
    .B(_16852_),
    .S(_05105_),
    .Z(_00777_));
 MUX2_X1 _30242_ (.A(_16981_),
    .B(_16853_),
    .S(_05105_),
    .Z(_00778_));
 MUX2_X1 _30243_ (.A(_16982_),
    .B(_16854_),
    .S(_05105_),
    .Z(_00779_));
 MUX2_X1 _30244_ (.A(_16983_),
    .B(_16855_),
    .S(_05105_),
    .Z(_00780_));
 MUX2_X1 _30245_ (.A(_16984_),
    .B(_16856_),
    .S(_05105_),
    .Z(_00781_));
 MUX2_X1 _30246_ (.A(_16986_),
    .B(_16858_),
    .S(_05105_),
    .Z(_00783_));
 BUF_X2 _30247_ (.A(_05104_),
    .Z(_05107_));
 MUX2_X1 _30248_ (.A(_16987_),
    .B(_16859_),
    .S(_05107_),
    .Z(_00784_));
 MUX2_X1 _30249_ (.A(_16988_),
    .B(_16860_),
    .S(_05107_),
    .Z(_00785_));
 MUX2_X1 _30250_ (.A(_16989_),
    .B(_16861_),
    .S(_05107_),
    .Z(_00786_));
 MUX2_X1 _30251_ (.A(_16990_),
    .B(_16862_),
    .S(_05107_),
    .Z(_00787_));
 MUX2_X1 _30252_ (.A(_16991_),
    .B(_16863_),
    .S(_05107_),
    .Z(_00788_));
 MUX2_X1 _30253_ (.A(_16992_),
    .B(_16864_),
    .S(_05107_),
    .Z(_00789_));
 MUX2_X1 _30254_ (.A(_16993_),
    .B(_16865_),
    .S(_05107_),
    .Z(_00790_));
 MUX2_X1 _30255_ (.A(_16994_),
    .B(_16866_),
    .S(_05107_),
    .Z(_00791_));
 MUX2_X1 _30256_ (.A(_16995_),
    .B(_16867_),
    .S(_05107_),
    .Z(_00792_));
 MUX2_X1 _30257_ (.A(_16997_),
    .B(_16869_),
    .S(_05107_),
    .Z(_00794_));
 BUF_X2 _30258_ (.A(_05104_),
    .Z(_05109_));
 MUX2_X1 _30259_ (.A(_16998_),
    .B(_16870_),
    .S(_05109_),
    .Z(_00795_));
 MUX2_X1 _30260_ (.A(_16999_),
    .B(_16871_),
    .S(_05109_),
    .Z(_00796_));
 MUX2_X1 _30261_ (.A(_17000_),
    .B(_16872_),
    .S(_05109_),
    .Z(_00797_));
 MUX2_X1 _30262_ (.A(_17001_),
    .B(_16873_),
    .S(_05109_),
    .Z(_00798_));
 MUX2_X1 _30263_ (.A(_17002_),
    .B(_16874_),
    .S(_05109_),
    .Z(_00799_));
 MUX2_X1 _30264_ (.A(_17003_),
    .B(_16875_),
    .S(_05109_),
    .Z(_00800_));
 MUX2_X1 _30265_ (.A(_17004_),
    .B(_16876_),
    .S(_05109_),
    .Z(_00801_));
 MUX2_X1 _30266_ (.A(_17005_),
    .B(_16877_),
    .S(_05109_),
    .Z(_00802_));
 MUX2_X1 _30267_ (.A(_17006_),
    .B(_16878_),
    .S(_05109_),
    .Z(_00803_));
 MUX2_X1 _30268_ (.A(_17008_),
    .B(_16880_),
    .S(_05109_),
    .Z(_00805_));
 BUF_X2 _30269_ (.A(_05104_),
    .Z(_05111_));
 MUX2_X1 _30270_ (.A(_17009_),
    .B(_16881_),
    .S(_05111_),
    .Z(_00806_));
 MUX2_X1 _30271_ (.A(_17010_),
    .B(_16882_),
    .S(_05111_),
    .Z(_00807_));
 MUX2_X1 _30272_ (.A(_17011_),
    .B(_16883_),
    .S(_05111_),
    .Z(_00808_));
 MUX2_X1 _30273_ (.A(_17012_),
    .B(_16884_),
    .S(_05111_),
    .Z(_00809_));
 MUX2_X1 _30274_ (.A(_17013_),
    .B(_16885_),
    .S(_05111_),
    .Z(_00810_));
 MUX2_X1 _30275_ (.A(_17014_),
    .B(_16886_),
    .S(_05111_),
    .Z(_00811_));
 MUX2_X1 _30276_ (.A(_17015_),
    .B(_16887_),
    .S(_05111_),
    .Z(_00812_));
 MUX2_X1 _30277_ (.A(_17016_),
    .B(_16888_),
    .S(_05111_),
    .Z(_00813_));
 MUX2_X1 _30278_ (.A(_17017_),
    .B(_16889_),
    .S(_05111_),
    .Z(_00814_));
 MUX2_X1 _30279_ (.A(_17019_),
    .B(_16891_),
    .S(_05111_),
    .Z(_00816_));
 BUF_X2 _30280_ (.A(_05104_),
    .Z(_05113_));
 MUX2_X1 _30281_ (.A(_17020_),
    .B(_16892_),
    .S(_05113_),
    .Z(_00817_));
 MUX2_X1 _30282_ (.A(_17021_),
    .B(_16893_),
    .S(_05113_),
    .Z(_00818_));
 MUX2_X1 _30283_ (.A(_17022_),
    .B(_16894_),
    .S(_05113_),
    .Z(_00819_));
 MUX2_X1 _30284_ (.A(_17023_),
    .B(_16895_),
    .S(_05113_),
    .Z(_00820_));
 MUX2_X1 _30285_ (.A(_17024_),
    .B(_16896_),
    .S(_05113_),
    .Z(_00821_));
 MUX2_X1 _30286_ (.A(_17025_),
    .B(_16897_),
    .S(_05113_),
    .Z(_00822_));
 MUX2_X1 _30287_ (.A(_17026_),
    .B(_16898_),
    .S(_05113_),
    .Z(_00823_));
 MUX2_X1 _30288_ (.A(_17027_),
    .B(_16899_),
    .S(_05113_),
    .Z(_00824_));
 MUX2_X1 _30289_ (.A(_17028_),
    .B(_16900_),
    .S(_05113_),
    .Z(_00825_));
 MUX2_X1 _30290_ (.A(_17030_),
    .B(_16902_),
    .S(_05113_),
    .Z(_00827_));
 BUF_X2 _30291_ (.A(_05104_),
    .Z(_05115_));
 MUX2_X1 _30292_ (.A(_17031_),
    .B(_16903_),
    .S(_05115_),
    .Z(_00828_));
 MUX2_X1 _30293_ (.A(_17032_),
    .B(_16904_),
    .S(_05115_),
    .Z(_00829_));
 MUX2_X1 _30294_ (.A(_17033_),
    .B(_16905_),
    .S(_05115_),
    .Z(_00830_));
 MUX2_X1 _30295_ (.A(_17034_),
    .B(_16906_),
    .S(_05115_),
    .Z(_00831_));
 MUX2_X1 _30296_ (.A(_17035_),
    .B(_16907_),
    .S(_05115_),
    .Z(_00832_));
 MUX2_X1 _30297_ (.A(_17036_),
    .B(_16908_),
    .S(_05115_),
    .Z(_00833_));
 MUX2_X1 _30298_ (.A(_17037_),
    .B(_16909_),
    .S(_05115_),
    .Z(_00834_));
 MUX2_X1 _30299_ (.A(_17038_),
    .B(_16910_),
    .S(_05115_),
    .Z(_00835_));
 MUX2_X1 _30300_ (.A(_17039_),
    .B(_16911_),
    .S(_05115_),
    .Z(_00836_));
 MUX2_X1 _30301_ (.A(_17041_),
    .B(_16913_),
    .S(_05115_),
    .Z(_00838_));
 BUF_X2 _30302_ (.A(_05104_),
    .Z(_05117_));
 MUX2_X1 _30303_ (.A(_17042_),
    .B(_16914_),
    .S(_05117_),
    .Z(_00839_));
 MUX2_X1 _30304_ (.A(_17043_),
    .B(_16915_),
    .S(_05117_),
    .Z(_00840_));
 MUX2_X1 _30305_ (.A(_17044_),
    .B(_16916_),
    .S(_05117_),
    .Z(_00841_));
 MUX2_X1 _30306_ (.A(_17045_),
    .B(_16917_),
    .S(_05117_),
    .Z(_00842_));
 MUX2_X1 _30307_ (.A(_17046_),
    .B(_16918_),
    .S(_05117_),
    .Z(_00843_));
 MUX2_X1 _30308_ (.A(_17047_),
    .B(_16919_),
    .S(_05117_),
    .Z(_00844_));
 MUX2_X1 _30309_ (.A(_17048_),
    .B(_16920_),
    .S(_05117_),
    .Z(_00845_));
 MUX2_X1 _30310_ (.A(_17049_),
    .B(_16921_),
    .S(_05117_),
    .Z(_00846_));
 MUX2_X1 _30311_ (.A(_17050_),
    .B(_16922_),
    .S(_05117_),
    .Z(_00847_));
 MUX2_X1 _30312_ (.A(_17052_),
    .B(_16924_),
    .S(_05117_),
    .Z(_00849_));
 BUF_X2 _30313_ (.A(_05104_),
    .Z(_05119_));
 MUX2_X1 _30314_ (.A(_17053_),
    .B(_16925_),
    .S(_05119_),
    .Z(_00850_));
 MUX2_X1 _30315_ (.A(_17054_),
    .B(_16926_),
    .S(_05119_),
    .Z(_00851_));
 MUX2_X1 _30316_ (.A(_17055_),
    .B(_16927_),
    .S(_05119_),
    .Z(_00852_));
 MUX2_X1 _30317_ (.A(_17056_),
    .B(_16928_),
    .S(_05119_),
    .Z(_00853_));
 MUX2_X1 _30318_ (.A(_17057_),
    .B(_16929_),
    .S(_05119_),
    .Z(_00854_));
 XOR2_X1 _30319_ (.A(_17099_),
    .B(_17058_),
    .Z(_05121_));
 BUF_X2 _30320_ (.A(_16680_),
    .Z(_05122_));
 AND2_X1 _30321_ (.A1(_05122_),
    .A2(_16679_),
    .ZN(_05123_));
 BUF_X2 _30322_ (.A(_05123_),
    .Z(_05124_));
 AND2_X2 _30323_ (.A1(_16681_),
    .A2(_16682_),
    .ZN(_05125_));
 AND2_X2 _30324_ (.A1(_05124_),
    .A2(_05125_),
    .ZN(_05127_));
 AND2_X1 _30325_ (.A1(_16684_),
    .A2(_16683_),
    .ZN(_05128_));
 CLKBUF_X2 _30326_ (.A(_05128_),
    .Z(_05129_));
 NOR2_X1 _30327_ (.A1(_16686_),
    .A2(_16685_),
    .ZN(_05130_));
 AND2_X1 _30328_ (.A1(_05129_),
    .A2(_05130_),
    .ZN(_05131_));
 AND2_X1 _30329_ (.A1(_05127_),
    .A2(_05131_),
    .ZN(_05132_));
 INV_X1 _30330_ (.A(_16682_),
    .ZN(_05133_));
 NOR2_X2 _30331_ (.A1(_05133_),
    .A2(_16681_),
    .ZN(_05134_));
 CLKBUF_X2 _30332_ (.A(_05134_),
    .Z(_05135_));
 NOR2_X2 _30333_ (.A1(_05122_),
    .A2(_16679_),
    .ZN(_05136_));
 BUF_X2 _30334_ (.A(_05136_),
    .Z(_05138_));
 AND3_X1 _30335_ (.A1(_05131_),
    .A2(_05135_),
    .A3(_05138_),
    .ZN(_05139_));
 INV_X2 _30336_ (.A(_16680_),
    .ZN(_05140_));
 AND2_X2 _30337_ (.A1(_05125_),
    .A2(_05140_),
    .ZN(_05141_));
 CLKBUF_X2 _30338_ (.A(_05141_),
    .Z(_05142_));
 BUF_X2 _30339_ (.A(_05131_),
    .Z(_05143_));
 AOI211_X1 _30340_ (.A(_05132_),
    .B(_05139_),
    .C1(_05142_),
    .C2(_05143_),
    .ZN(_05144_));
 NOR2_X2 _30341_ (.A1(_05140_),
    .A2(_16679_),
    .ZN(_05145_));
 CLKBUF_X2 _30342_ (.A(_05145_),
    .Z(_05146_));
 INV_X1 _30343_ (.A(_16681_),
    .ZN(_05147_));
 NOR2_X2 _30344_ (.A1(_05147_),
    .A2(_16682_),
    .ZN(_05149_));
 BUF_X2 _30345_ (.A(_05149_),
    .Z(_05150_));
 BUF_X2 _30346_ (.A(_05129_),
    .Z(_05151_));
 BUF_X2 _30347_ (.A(_05130_),
    .Z(_05152_));
 NAND4_X1 _30348_ (.A1(_05146_),
    .A2(_05150_),
    .A3(_05151_),
    .A4(_05152_),
    .ZN(_05153_));
 INV_X1 _30349_ (.A(_05131_),
    .ZN(_05154_));
 INV_X1 _30350_ (.A(_05136_),
    .ZN(_05155_));
 NOR2_X1 _30351_ (.A1(_16681_),
    .A2(_16682_),
    .ZN(_05156_));
 CLKBUF_X2 _30352_ (.A(_05156_),
    .Z(_05157_));
 NAND2_X1 _30353_ (.A1(_05155_),
    .A2(_05157_),
    .ZN(_05158_));
 OAI211_X1 _30354_ (.A(_05144_),
    .B(_05153_),
    .C1(_05154_),
    .C2(_05158_),
    .ZN(_05160_));
 NOR2_X1 _30355_ (.A1(_16684_),
    .A2(_16683_),
    .ZN(_05161_));
 AND2_X1 _30356_ (.A1(_05161_),
    .A2(_05130_),
    .ZN(_05162_));
 CLKBUF_X2 _30357_ (.A(_05162_),
    .Z(_05163_));
 BUF_X2 _30358_ (.A(_05122_),
    .Z(_05164_));
 CLKBUF_X2 _30359_ (.A(_16679_),
    .Z(_05165_));
 BUF_X2 _30360_ (.A(_05165_),
    .Z(_05166_));
 OAI211_X1 _30361_ (.A(_05163_),
    .B(_05150_),
    .C1(_05164_),
    .C2(_05166_),
    .ZN(_05167_));
 CLKBUF_X2 _30362_ (.A(_05135_),
    .Z(_05168_));
 OAI211_X1 _30363_ (.A(_05163_),
    .B(_05168_),
    .C1(_05164_),
    .C2(_05166_),
    .ZN(_05169_));
 CLKBUF_X2 _30364_ (.A(_05125_),
    .Z(_05171_));
 INV_X2 _30365_ (.A(_16679_),
    .ZN(_05172_));
 NOR2_X2 _30366_ (.A1(_05172_),
    .A2(_05122_),
    .ZN(_05173_));
 OAI211_X1 _30367_ (.A(_05163_),
    .B(_05171_),
    .C1(_05146_),
    .C2(_05173_),
    .ZN(_05174_));
 CLKBUF_X2 _30368_ (.A(_05163_),
    .Z(_05175_));
 AND2_X1 _30369_ (.A1(_05157_),
    .A2(_05122_),
    .ZN(_05176_));
 BUF_X2 _30370_ (.A(_05176_),
    .Z(_05177_));
 NAND2_X1 _30371_ (.A1(_05175_),
    .A2(_05177_),
    .ZN(_05178_));
 NAND4_X1 _30372_ (.A1(_05167_),
    .A2(_05169_),
    .A3(_05174_),
    .A4(_05178_),
    .ZN(_05179_));
 NOR3_X2 _30373_ (.A1(_05145_),
    .A2(_16681_),
    .A3(_05133_),
    .ZN(_05180_));
 INV_X1 _30374_ (.A(_05173_),
    .ZN(_05182_));
 AND2_X1 _30375_ (.A1(_05180_),
    .A2(_05182_),
    .ZN(_05183_));
 INV_X1 _30376_ (.A(_16683_),
    .ZN(_05184_));
 NOR2_X1 _30377_ (.A1(_05184_),
    .A2(_16684_),
    .ZN(_05185_));
 AND2_X1 _30378_ (.A1(_05185_),
    .A2(_05130_),
    .ZN(_05186_));
 BUF_X2 _30379_ (.A(_05186_),
    .Z(_05187_));
 NAND2_X1 _30380_ (.A1(_05183_),
    .A2(_05187_),
    .ZN(_05188_));
 NAND2_X1 _30381_ (.A1(_05187_),
    .A2(_05177_),
    .ZN(_05189_));
 INV_X2 _30382_ (.A(_05124_),
    .ZN(_05190_));
 NAND2_X1 _30383_ (.A1(_05190_),
    .A2(_05149_),
    .ZN(_05191_));
 NOR2_X1 _30384_ (.A1(_05191_),
    .A2(_05138_),
    .ZN(_05193_));
 INV_X1 _30385_ (.A(_05193_),
    .ZN(_05194_));
 INV_X1 _30386_ (.A(_05186_),
    .ZN(_05195_));
 OAI211_X1 _30387_ (.A(_05188_),
    .B(_05189_),
    .C1(_05194_),
    .C2(_05195_),
    .ZN(_05196_));
 AND2_X1 _30388_ (.A1(_05184_),
    .A2(_16684_),
    .ZN(_05197_));
 AND2_X1 _30389_ (.A1(_05197_),
    .A2(_05130_),
    .ZN(_05198_));
 BUF_X2 _30390_ (.A(_05198_),
    .Z(_05199_));
 BUF_X2 _30391_ (.A(_05157_),
    .Z(_05200_));
 NOR3_X1 _30392_ (.A1(_05136_),
    .A2(_05147_),
    .A3(_16682_),
    .ZN(_05201_));
 OAI211_X1 _30393_ (.A(_05199_),
    .B(_05190_),
    .C1(_05200_),
    .C2(_05201_),
    .ZN(_05202_));
 AND2_X1 _30394_ (.A1(_05155_),
    .A2(_05134_),
    .ZN(_05204_));
 NAND2_X1 _30395_ (.A1(_05198_),
    .A2(_05204_),
    .ZN(_05205_));
 CLKBUF_X2 _30396_ (.A(_05197_),
    .Z(_05206_));
 AND2_X1 _30397_ (.A1(_05125_),
    .A2(_05122_),
    .ZN(_05207_));
 AND2_X1 _30398_ (.A1(_05125_),
    .A2(_05136_),
    .ZN(_05208_));
 BUF_X2 _30399_ (.A(_05208_),
    .Z(_05209_));
 OAI211_X1 _30400_ (.A(_05206_),
    .B(_05152_),
    .C1(_05207_),
    .C2(_05209_),
    .ZN(_05210_));
 NAND3_X1 _30401_ (.A1(_05202_),
    .A2(_05205_),
    .A3(_05210_),
    .ZN(_05211_));
 NOR4_X1 _30402_ (.A1(_05160_),
    .A2(_05179_),
    .A3(_05196_),
    .A4(_05211_),
    .ZN(_05212_));
 AND2_X2 _30403_ (.A1(_05145_),
    .A2(_05156_),
    .ZN(_05213_));
 CLKBUF_X2 _30404_ (.A(_05185_),
    .Z(_05215_));
 AND2_X1 _30405_ (.A1(_16686_),
    .A2(_16685_),
    .ZN(_05216_));
 AND2_X2 _30406_ (.A1(_05215_),
    .A2(_05216_),
    .ZN(_05217_));
 NAND2_X1 _30407_ (.A1(_05213_),
    .A2(_05217_),
    .ZN(_05218_));
 AND2_X2 _30408_ (.A1(_05173_),
    .A2(_05149_),
    .ZN(_05219_));
 BUF_X2 _30409_ (.A(_05217_),
    .Z(_05220_));
 NAND2_X1 _30410_ (.A1(_05219_),
    .A2(_05220_),
    .ZN(_05221_));
 NAND2_X1 _30411_ (.A1(_05218_),
    .A2(_05221_),
    .ZN(_05222_));
 AND2_X1 _30412_ (.A1(_05216_),
    .A2(_05161_),
    .ZN(_05223_));
 AND3_X1 _30413_ (.A1(_05223_),
    .A2(_05165_),
    .A3(_05134_),
    .ZN(_05224_));
 AND2_X1 _30414_ (.A1(_05141_),
    .A2(_05223_),
    .ZN(_05226_));
 CLKBUF_X2 _30415_ (.A(_05161_),
    .Z(_05227_));
 AND4_X1 _30416_ (.A1(_05145_),
    .A2(_05125_),
    .A3(_05227_),
    .A4(_05216_),
    .ZN(_05228_));
 OR3_X1 _30417_ (.A1(_05224_),
    .A2(_05226_),
    .A3(_05228_),
    .ZN(_05229_));
 AND2_X1 _30418_ (.A1(_05134_),
    .A2(_05140_),
    .ZN(_05230_));
 NAND2_X1 _30419_ (.A1(_05230_),
    .A2(_05217_),
    .ZN(_05231_));
 AND2_X2 _30420_ (.A1(_05134_),
    .A2(_05122_),
    .ZN(_05232_));
 NAND2_X1 _30421_ (.A1(_05232_),
    .A2(_05217_),
    .ZN(_05233_));
 AND2_X1 _30422_ (.A1(_05145_),
    .A2(_05125_),
    .ZN(_05234_));
 BUF_X2 _30423_ (.A(_05234_),
    .Z(_05235_));
 AND2_X2 _30424_ (.A1(_05173_),
    .A2(_05125_),
    .ZN(_05237_));
 NOR2_X1 _30425_ (.A1(_05235_),
    .A2(_05237_),
    .ZN(_05238_));
 INV_X1 _30426_ (.A(_05217_),
    .ZN(_05239_));
 OAI211_X1 _30427_ (.A(_05231_),
    .B(_05233_),
    .C1(_05238_),
    .C2(_05239_),
    .ZN(_05240_));
 AND4_X1 _30428_ (.A1(_05145_),
    .A2(_05157_),
    .A3(_05227_),
    .A4(_05216_),
    .ZN(_05241_));
 OR4_X1 _30429_ (.A1(_05222_),
    .A2(_05229_),
    .A3(_05240_),
    .A4(_05241_),
    .ZN(_05242_));
 AND2_X2 _30430_ (.A1(_05197_),
    .A2(_05216_),
    .ZN(_05243_));
 BUF_X2 _30431_ (.A(_05243_),
    .Z(_05244_));
 AND2_X1 _30432_ (.A1(_05124_),
    .A2(_05156_),
    .ZN(_05245_));
 INV_X1 _30433_ (.A(_05245_),
    .ZN(_05246_));
 AND2_X2 _30434_ (.A1(_05136_),
    .A2(_05156_),
    .ZN(_05248_));
 INV_X1 _30435_ (.A(_05248_),
    .ZN(_05249_));
 NAND2_X2 _30436_ (.A1(_05246_),
    .A2(_05249_),
    .ZN(_05250_));
 AND2_X1 _30437_ (.A1(_05149_),
    .A2(_05140_),
    .ZN(_05251_));
 BUF_X2 _30438_ (.A(_05251_),
    .Z(_05252_));
 OAI21_X1 _30439_ (.A(_05244_),
    .B1(_05250_),
    .B2(_05252_),
    .ZN(_05253_));
 NAND3_X1 _30440_ (.A1(_05243_),
    .A2(_05135_),
    .A3(_05182_),
    .ZN(_05254_));
 INV_X1 _30441_ (.A(_05243_),
    .ZN(_05255_));
 AND2_X1 _30442_ (.A1(_05125_),
    .A2(_16679_),
    .ZN(_05256_));
 INV_X1 _30443_ (.A(_05256_),
    .ZN(_05257_));
 OAI211_X1 _30444_ (.A(_05253_),
    .B(_05254_),
    .C1(_05255_),
    .C2(_05257_),
    .ZN(_05259_));
 AND2_X1 _30445_ (.A1(_05173_),
    .A2(_05157_),
    .ZN(_05260_));
 BUF_X2 _30446_ (.A(_05260_),
    .Z(_05261_));
 AND2_X2 _30447_ (.A1(_05129_),
    .A2(_05216_),
    .ZN(_05262_));
 BUF_X2 _30448_ (.A(_05262_),
    .Z(_05263_));
 NAND2_X1 _30449_ (.A1(_05261_),
    .A2(_05263_),
    .ZN(_05264_));
 AND2_X1 _30450_ (.A1(_05149_),
    .A2(_05136_),
    .ZN(_05265_));
 NAND2_X1 _30451_ (.A1(_05265_),
    .A2(_05262_),
    .ZN(_05266_));
 CLKBUF_X2 _30452_ (.A(_05216_),
    .Z(_05267_));
 NAND3_X1 _30453_ (.A1(_05177_),
    .A2(_05151_),
    .A3(_05267_),
    .ZN(_05268_));
 NAND3_X1 _30454_ (.A1(_05264_),
    .A2(_05266_),
    .A3(_05268_),
    .ZN(_05270_));
 NAND2_X1 _30455_ (.A1(_05232_),
    .A2(_05262_),
    .ZN(_05271_));
 NAND3_X1 _30456_ (.A1(_05262_),
    .A2(_05146_),
    .A3(_05171_),
    .ZN(_05272_));
 INV_X1 _30457_ (.A(_05230_),
    .ZN(_05273_));
 INV_X1 _30458_ (.A(_05262_),
    .ZN(_05274_));
 OAI211_X1 _30459_ (.A(_05271_),
    .B(_05272_),
    .C1(_05273_),
    .C2(_05274_),
    .ZN(_05275_));
 NOR4_X1 _30460_ (.A1(_05242_),
    .A2(_05259_),
    .A3(_05270_),
    .A4(_05275_),
    .ZN(_05276_));
 INV_X1 _30461_ (.A(_16686_),
    .ZN(_05277_));
 AND2_X1 _30462_ (.A1(_05277_),
    .A2(_16685_),
    .ZN(_05278_));
 AND2_X1 _30463_ (.A1(_05278_),
    .A2(_05161_),
    .ZN(_05279_));
 BUF_X2 _30464_ (.A(_05279_),
    .Z(_05281_));
 OAI21_X1 _30465_ (.A(_05281_),
    .B1(_05235_),
    .B2(_05142_),
    .ZN(_05282_));
 AND2_X1 _30466_ (.A1(_05156_),
    .A2(_05140_),
    .ZN(_05283_));
 BUF_X2 _30467_ (.A(_05283_),
    .Z(_05284_));
 OAI21_X1 _30468_ (.A(_05281_),
    .B1(_05265_),
    .B2(_05284_),
    .ZN(_05285_));
 CLKBUF_X2 _30469_ (.A(_05278_),
    .Z(_05286_));
 NAND4_X1 _30470_ (.A1(_05286_),
    .A2(_05135_),
    .A3(_05165_),
    .A4(_05227_),
    .ZN(_05287_));
 AND3_X1 _30471_ (.A1(_05282_),
    .A2(_05285_),
    .A3(_05287_),
    .ZN(_05288_));
 AND2_X1 _30472_ (.A1(_05197_),
    .A2(_05286_),
    .ZN(_05289_));
 AND2_X1 _30473_ (.A1(_05289_),
    .A2(_05235_),
    .ZN(_05290_));
 INV_X1 _30474_ (.A(_05289_),
    .ZN(_05292_));
 AND2_X1 _30475_ (.A1(_05156_),
    .A2(_05165_),
    .ZN(_05293_));
 INV_X1 _30476_ (.A(_05293_),
    .ZN(_05294_));
 INV_X1 _30477_ (.A(_05150_),
    .ZN(_05295_));
 AOI21_X1 _30478_ (.A(_05292_),
    .B1(_05294_),
    .B2(_05295_),
    .ZN(_05296_));
 BUF_X2 _30479_ (.A(_05289_),
    .Z(_05297_));
 AOI211_X1 _30480_ (.A(_05290_),
    .B(_05296_),
    .C1(_05297_),
    .C2(_05180_),
    .ZN(_05298_));
 AND2_X1 _30481_ (.A1(_05286_),
    .A2(_05215_),
    .ZN(_05299_));
 AND2_X1 _30482_ (.A1(_05149_),
    .A2(_05122_),
    .ZN(_05300_));
 CLKBUF_X2 _30483_ (.A(_05300_),
    .Z(_05301_));
 NAND2_X1 _30484_ (.A1(_05299_),
    .A2(_05301_),
    .ZN(_05303_));
 AND2_X1 _30485_ (.A1(_05299_),
    .A2(_05245_),
    .ZN(_05304_));
 INV_X1 _30486_ (.A(_05304_),
    .ZN(_05305_));
 AND2_X1 _30487_ (.A1(_05135_),
    .A2(_05165_),
    .ZN(_05306_));
 OAI21_X1 _30488_ (.A(_05299_),
    .B1(_05306_),
    .B2(_05127_),
    .ZN(_05307_));
 NAND2_X1 _30489_ (.A1(_05299_),
    .A2(_05284_),
    .ZN(_05308_));
 AND4_X1 _30490_ (.A1(_05303_),
    .A2(_05305_),
    .A3(_05307_),
    .A4(_05308_),
    .ZN(_05309_));
 AND2_X1 _30491_ (.A1(_05278_),
    .A2(_05129_),
    .ZN(_05310_));
 CLKBUF_X2 _30492_ (.A(_05310_),
    .Z(_05311_));
 BUF_X2 _30493_ (.A(_05245_),
    .Z(_05312_));
 NAND2_X1 _30494_ (.A1(_05311_),
    .A2(_05312_),
    .ZN(_05314_));
 AND2_X1 _30495_ (.A1(_05134_),
    .A2(_05123_),
    .ZN(_05315_));
 BUF_X2 _30496_ (.A(_05315_),
    .Z(_05316_));
 OAI21_X1 _30497_ (.A(_05310_),
    .B1(_05234_),
    .B2(_05316_),
    .ZN(_05317_));
 NAND3_X1 _30498_ (.A1(_05310_),
    .A2(_05165_),
    .A3(_05141_),
    .ZN(_05318_));
 AND2_X1 _30499_ (.A1(_05317_),
    .A2(_05318_),
    .ZN(_05319_));
 AND2_X1 _30500_ (.A1(_05149_),
    .A2(_05165_),
    .ZN(_05320_));
 NAND3_X1 _30501_ (.A1(_05320_),
    .A2(_05286_),
    .A3(_05129_),
    .ZN(_05321_));
 NAND3_X1 _30502_ (.A1(_05284_),
    .A2(_05286_),
    .A3(_05129_),
    .ZN(_05322_));
 AND4_X1 _30503_ (.A1(_05314_),
    .A2(_05319_),
    .A3(_05321_),
    .A4(_05322_),
    .ZN(_05323_));
 AND4_X1 _30504_ (.A1(_05288_),
    .A2(_05298_),
    .A3(_05309_),
    .A4(_05323_),
    .ZN(_05325_));
 NOR2_X1 _30505_ (.A1(_05277_),
    .A2(_16685_),
    .ZN(_05326_));
 CLKBUF_X2 _30506_ (.A(_05326_),
    .Z(_05327_));
 AND2_X1 _30507_ (.A1(_05215_),
    .A2(_05327_),
    .ZN(_05328_));
 CLKBUF_X2 _30508_ (.A(_05328_),
    .Z(_05329_));
 INV_X1 _30509_ (.A(_05157_),
    .ZN(_05330_));
 NOR3_X1 _30510_ (.A1(_05330_),
    .A2(_05124_),
    .A3(_05138_),
    .ZN(_05331_));
 BUF_X2 _30511_ (.A(_05207_),
    .Z(_05332_));
 OAI21_X1 _30512_ (.A(_05329_),
    .B1(_05331_),
    .B2(_05332_),
    .ZN(_05333_));
 OAI211_X1 _30513_ (.A(_05327_),
    .B(_05197_),
    .C1(_05127_),
    .C2(_05141_),
    .ZN(_05334_));
 NAND4_X1 _30514_ (.A1(_05197_),
    .A2(_05135_),
    .A3(_05173_),
    .A4(_05327_),
    .ZN(_05336_));
 INV_X1 _30515_ (.A(_05265_),
    .ZN(_05337_));
 AND2_X1 _30516_ (.A1(_05197_),
    .A2(_05327_),
    .ZN(_05338_));
 INV_X1 _30517_ (.A(_05338_),
    .ZN(_05339_));
 OAI211_X1 _30518_ (.A(_05334_),
    .B(_05336_),
    .C1(_05337_),
    .C2(_05339_),
    .ZN(_05340_));
 AND2_X1 _30519_ (.A1(_05326_),
    .A2(_05129_),
    .ZN(_05341_));
 INV_X2 _30520_ (.A(_05341_),
    .ZN(_05342_));
 INV_X1 _30521_ (.A(_05145_),
    .ZN(_05343_));
 NAND2_X1 _30522_ (.A1(_05343_),
    .A2(_05149_),
    .ZN(_05344_));
 NOR2_X1 _30523_ (.A1(_05342_),
    .A2(_05344_),
    .ZN(_05345_));
 CLKBUF_X2 _30524_ (.A(_05341_),
    .Z(_05347_));
 NOR2_X1 _30525_ (.A1(_05330_),
    .A2(_05173_),
    .ZN(_05348_));
 AND2_X1 _30526_ (.A1(_05347_),
    .A2(_05348_),
    .ZN(_05349_));
 AND3_X1 _30527_ (.A1(_05209_),
    .A2(_05129_),
    .A3(_05327_),
    .ZN(_05350_));
 NOR4_X1 _30528_ (.A1(_05340_),
    .A2(_05345_),
    .A3(_05349_),
    .A4(_05350_),
    .ZN(_05351_));
 AND2_X1 _30529_ (.A1(_05327_),
    .A2(_05161_),
    .ZN(_05352_));
 CLKBUF_X2 _30530_ (.A(_05352_),
    .Z(_05353_));
 NAND2_X1 _30531_ (.A1(_05353_),
    .A2(_05251_),
    .ZN(_05354_));
 NAND4_X1 _30532_ (.A1(_05150_),
    .A2(_05327_),
    .A3(_05124_),
    .A4(_05227_),
    .ZN(_05355_));
 NAND2_X1 _30533_ (.A1(_05354_),
    .A2(_05355_),
    .ZN(_05356_));
 BUF_X2 _30534_ (.A(_05353_),
    .Z(_05358_));
 AND2_X1 _30535_ (.A1(_05200_),
    .A2(_05172_),
    .ZN(_05359_));
 AOI21_X1 _30536_ (.A(_05356_),
    .B1(_05358_),
    .B2(_05359_),
    .ZN(_05360_));
 OAI21_X1 _30537_ (.A(_05125_),
    .B1(_05122_),
    .B2(_05165_),
    .ZN(_05361_));
 INV_X1 _30538_ (.A(_05361_),
    .ZN(_05362_));
 OAI21_X1 _30539_ (.A(_05358_),
    .B1(_05362_),
    .B2(_05306_),
    .ZN(_05363_));
 AND4_X1 _30540_ (.A1(_05333_),
    .A2(_05351_),
    .A3(_05360_),
    .A4(_05363_),
    .ZN(_05364_));
 AND4_X1 _30541_ (.A1(_05212_),
    .A2(_05276_),
    .A3(_05325_),
    .A4(_05364_),
    .ZN(_05365_));
 AND2_X1 _30542_ (.A1(_05248_),
    .A2(_05163_),
    .ZN(_05366_));
 INV_X1 _30543_ (.A(_05366_),
    .ZN(_05367_));
 NAND2_X2 _30544_ (.A1(_05365_),
    .A2(_05367_),
    .ZN(_05369_));
 AND2_X1 _30545_ (.A1(_05135_),
    .A2(_05173_),
    .ZN(_05370_));
 AND2_X1 _30546_ (.A1(_05370_),
    .A2(_05262_),
    .ZN(_05371_));
 INV_X1 _30547_ (.A(_05371_),
    .ZN(_05372_));
 NAND2_X1 _30548_ (.A1(_05289_),
    .A2(_05370_),
    .ZN(_05373_));
 NAND3_X1 _30549_ (.A1(_05262_),
    .A2(_05190_),
    .A3(_05200_),
    .ZN(_05374_));
 NAND2_X1 _30550_ (.A1(_05198_),
    .A2(_05237_),
    .ZN(_05375_));
 NAND4_X1 _30551_ (.A1(_05372_),
    .A2(_05373_),
    .A3(_05374_),
    .A4(_05375_),
    .ZN(_05376_));
 NAND3_X1 _30552_ (.A1(_05235_),
    .A2(_05327_),
    .A3(_05206_),
    .ZN(_05377_));
 INV_X1 _30553_ (.A(_05237_),
    .ZN(_05378_));
 BUF_X2 _30554_ (.A(_05223_),
    .Z(_05380_));
 INV_X1 _30555_ (.A(_05380_),
    .ZN(_05381_));
 OAI221_X1 _30556_ (.A(_05377_),
    .B1(_05378_),
    .B2(_05381_),
    .C1(_05339_),
    .C2(_05249_),
    .ZN(_05382_));
 AND2_X1 _30557_ (.A1(_05134_),
    .A2(_05145_),
    .ZN(_05383_));
 BUF_X2 _30558_ (.A(_05383_),
    .Z(_05384_));
 AOI22_X1 _30559_ (.A1(_05384_),
    .A2(_05338_),
    .B1(_05219_),
    .B2(_05353_),
    .ZN(_05385_));
 NAND2_X1 _30560_ (.A1(_05316_),
    .A2(_05217_),
    .ZN(_05386_));
 NAND4_X1 _30561_ (.A1(_05206_),
    .A2(_05133_),
    .A3(_05146_),
    .A4(_05267_),
    .ZN(_05387_));
 NAND3_X1 _30562_ (.A1(_05385_),
    .A2(_05386_),
    .A3(_05387_),
    .ZN(_05388_));
 AND2_X2 _30563_ (.A1(_05149_),
    .A2(_05124_),
    .ZN(_05389_));
 NAND2_X1 _30564_ (.A1(_05289_),
    .A2(_05389_),
    .ZN(_05391_));
 NAND2_X1 _30565_ (.A1(_05310_),
    .A2(_05293_),
    .ZN(_05392_));
 INV_X1 _30566_ (.A(_05310_),
    .ZN(_05393_));
 INV_X1 _30567_ (.A(_05389_),
    .ZN(_05394_));
 OAI211_X1 _30568_ (.A(_05391_),
    .B(_05392_),
    .C1(_05393_),
    .C2(_05394_),
    .ZN(_05395_));
 NOR4_X1 _30569_ (.A1(_05376_),
    .A2(_05382_),
    .A3(_05388_),
    .A4(_05395_),
    .ZN(_05396_));
 NAND2_X1 _30570_ (.A1(_05289_),
    .A2(_05200_),
    .ZN(_05397_));
 AND2_X1 _30571_ (.A1(_05187_),
    .A2(_05141_),
    .ZN(_05398_));
 INV_X1 _30572_ (.A(_05127_),
    .ZN(_05399_));
 INV_X1 _30573_ (.A(_05213_),
    .ZN(_05400_));
 AOI21_X1 _30574_ (.A(_05195_),
    .B1(_05399_),
    .B2(_05400_),
    .ZN(_05402_));
 AOI211_X1 _30575_ (.A(_05398_),
    .B(_05402_),
    .C1(_05232_),
    .C2(_05187_),
    .ZN(_05403_));
 NAND2_X1 _30576_ (.A1(_05142_),
    .A2(_05163_),
    .ZN(_05404_));
 AOI22_X1 _30577_ (.A1(_05207_),
    .A2(_05289_),
    .B1(_05311_),
    .B2(_05251_),
    .ZN(_05405_));
 AND4_X1 _30578_ (.A1(_05397_),
    .A2(_05403_),
    .A3(_05404_),
    .A4(_05405_),
    .ZN(_05406_));
 NOR2_X1 _30579_ (.A1(_05344_),
    .A2(_05173_),
    .ZN(_05407_));
 OAI21_X1 _30580_ (.A(_05163_),
    .B1(_05407_),
    .B2(_05235_),
    .ZN(_05408_));
 OAI21_X1 _30581_ (.A(_05380_),
    .B1(_05201_),
    .B2(_05248_),
    .ZN(_05409_));
 AND3_X1 _30582_ (.A1(_05254_),
    .A2(_05205_),
    .A3(_05409_),
    .ZN(_05410_));
 AND2_X1 _30583_ (.A1(_05310_),
    .A2(_05362_),
    .ZN(_05411_));
 INV_X1 _30584_ (.A(_05411_),
    .ZN(_05413_));
 AND2_X1 _30585_ (.A1(_05171_),
    .A2(_05172_),
    .ZN(_05414_));
 OAI21_X1 _30586_ (.A(_05131_),
    .B1(_05232_),
    .B2(_05414_),
    .ZN(_05415_));
 AND4_X1 _30587_ (.A1(_05408_),
    .A2(_05410_),
    .A3(_05413_),
    .A4(_05415_),
    .ZN(_05416_));
 NAND2_X1 _30588_ (.A1(_05234_),
    .A2(_05347_),
    .ZN(_05417_));
 NAND2_X1 _30589_ (.A1(_05232_),
    .A2(_05341_),
    .ZN(_05418_));
 NAND2_X1 _30590_ (.A1(_05417_),
    .A2(_05418_),
    .ZN(_05419_));
 AND3_X1 _30591_ (.A1(_05217_),
    .A2(_05343_),
    .A3(_05171_),
    .ZN(_05420_));
 OR3_X1 _30592_ (.A1(_05419_),
    .A2(_05345_),
    .A3(_05420_),
    .ZN(_05421_));
 AND2_X1 _30593_ (.A1(_05310_),
    .A2(_05383_),
    .ZN(_05422_));
 AND2_X1 _30594_ (.A1(_05311_),
    .A2(_05230_),
    .ZN(_05424_));
 NAND3_X1 _30595_ (.A1(_05283_),
    .A2(_05206_),
    .A3(_05152_),
    .ZN(_05425_));
 NAND4_X1 _30596_ (.A1(_05197_),
    .A2(_05146_),
    .A3(_05157_),
    .A4(_05152_),
    .ZN(_05426_));
 NAND2_X1 _30597_ (.A1(_05425_),
    .A2(_05426_),
    .ZN(_05427_));
 NOR4_X1 _30598_ (.A1(_05421_),
    .A2(_05422_),
    .A3(_05424_),
    .A4(_05427_),
    .ZN(_05428_));
 AND4_X1 _30599_ (.A1(_05396_),
    .A2(_05406_),
    .A3(_05416_),
    .A4(_05428_),
    .ZN(_05429_));
 AND2_X1 _30600_ (.A1(_05204_),
    .A2(_05190_),
    .ZN(_05430_));
 AND2_X1 _30601_ (.A1(_05430_),
    .A2(_05328_),
    .ZN(_05431_));
 INV_X1 _30602_ (.A(_05328_),
    .ZN(_05432_));
 INV_X1 _30603_ (.A(_05301_),
    .ZN(_05433_));
 AOI21_X1 _30604_ (.A(_05432_),
    .B1(_05294_),
    .B2(_05433_),
    .ZN(_05435_));
 INV_X1 _30605_ (.A(_05208_),
    .ZN(_05436_));
 AOI21_X1 _30606_ (.A(_05432_),
    .B1(_05399_),
    .B2(_05436_),
    .ZN(_05437_));
 CLKBUF_X2 _30607_ (.A(_05327_),
    .Z(_05438_));
 AND3_X1 _30608_ (.A1(_05141_),
    .A2(_05438_),
    .A3(_05206_),
    .ZN(_05439_));
 NOR4_X1 _30609_ (.A1(_05431_),
    .A2(_05435_),
    .A3(_05437_),
    .A4(_05439_),
    .ZN(_05440_));
 BUF_X2 _30610_ (.A(_05299_),
    .Z(_05441_));
 OAI21_X1 _30611_ (.A(_05441_),
    .B1(_05430_),
    .B2(_05127_),
    .ZN(_05442_));
 NAND4_X1 _30612_ (.A1(_05286_),
    .A2(_05215_),
    .A3(_05165_),
    .A4(_05157_),
    .ZN(_05443_));
 AND2_X1 _30613_ (.A1(_05145_),
    .A2(_05149_),
    .ZN(_05444_));
 BUF_X2 _30614_ (.A(_05444_),
    .Z(_05446_));
 OAI21_X1 _30615_ (.A(_05299_),
    .B1(_05219_),
    .B2(_05446_),
    .ZN(_05447_));
 NAND3_X1 _30616_ (.A1(_05442_),
    .A2(_05443_),
    .A3(_05447_),
    .ZN(_05448_));
 INV_X1 _30617_ (.A(_05283_),
    .ZN(_05449_));
 OAI22_X1 _30618_ (.A1(_05339_),
    .A2(_05273_),
    .B1(_05342_),
    .B2(_05449_),
    .ZN(_05450_));
 INV_X1 _30619_ (.A(_05281_),
    .ZN(_05451_));
 INV_X1 _30620_ (.A(_05260_),
    .ZN(_05452_));
 AOI21_X1 _30621_ (.A(_05451_),
    .B1(_05452_),
    .B2(_05394_),
    .ZN(_05453_));
 INV_X1 _30622_ (.A(_05232_),
    .ZN(_05454_));
 AOI21_X1 _30623_ (.A(_05451_),
    .B1(_05454_),
    .B2(_05257_),
    .ZN(_05455_));
 NOR4_X1 _30624_ (.A1(_05448_),
    .A2(_05450_),
    .A3(_05453_),
    .A4(_05455_),
    .ZN(_05457_));
 NAND2_X1 _30625_ (.A1(_05399_),
    .A2(_05436_),
    .ZN(_05458_));
 NAND2_X1 _30626_ (.A1(_05458_),
    .A2(_05243_),
    .ZN(_05459_));
 NAND2_X1 _30627_ (.A1(_05243_),
    .A2(_05284_),
    .ZN(_05460_));
 NAND2_X1 _30628_ (.A1(_05243_),
    .A2(_05320_),
    .ZN(_05461_));
 BUF_X2 _30629_ (.A(_05230_),
    .Z(_05462_));
 OAI21_X1 _30630_ (.A(_05462_),
    .B1(_05353_),
    .B2(_05380_),
    .ZN(_05463_));
 NAND4_X1 _30631_ (.A1(_05459_),
    .A2(_05460_),
    .A3(_05461_),
    .A4(_05463_),
    .ZN(_05464_));
 NAND2_X1 _30632_ (.A1(_05250_),
    .A2(_05353_),
    .ZN(_05465_));
 AND2_X1 _30633_ (.A1(_05207_),
    .A2(_05223_),
    .ZN(_05466_));
 INV_X1 _30634_ (.A(_05466_),
    .ZN(_05468_));
 NAND2_X1 _30635_ (.A1(_05446_),
    .A2(_05217_),
    .ZN(_05469_));
 NAND4_X1 _30636_ (.A1(_05465_),
    .A2(_05468_),
    .A3(_05218_),
    .A4(_05469_),
    .ZN(_05470_));
 AND2_X1 _30637_ (.A1(_05198_),
    .A2(_05300_),
    .ZN(_05471_));
 NAND2_X1 _30638_ (.A1(_05187_),
    .A2(_05230_),
    .ZN(_05472_));
 NAND2_X1 _30639_ (.A1(_05187_),
    .A2(_05283_),
    .ZN(_05473_));
 NAND2_X1 _30640_ (.A1(_05472_),
    .A2(_05473_),
    .ZN(_05474_));
 NOR4_X1 _30641_ (.A1(_05464_),
    .A2(_05470_),
    .A3(_05471_),
    .A4(_05474_),
    .ZN(_05475_));
 AND2_X1 _30642_ (.A1(_05407_),
    .A2(_05187_),
    .ZN(_05476_));
 INV_X1 _30643_ (.A(_05251_),
    .ZN(_05477_));
 OAI22_X1 _30644_ (.A1(_05477_),
    .A2(_05274_),
    .B1(_05154_),
    .B2(_05294_),
    .ZN(_05479_));
 AND2_X1 _30645_ (.A1(_05320_),
    .A2(_05131_),
    .ZN(_05480_));
 AND2_X1 _30646_ (.A1(_05262_),
    .A2(_05414_),
    .ZN(_05481_));
 NOR4_X1 _30647_ (.A1(_05476_),
    .A2(_05479_),
    .A3(_05480_),
    .A4(_05481_),
    .ZN(_05482_));
 AND4_X1 _30648_ (.A1(_05440_),
    .A2(_05457_),
    .A3(_05475_),
    .A4(_05482_),
    .ZN(_05483_));
 AND2_X2 _30649_ (.A1(_05429_),
    .A2(_05483_),
    .ZN(_05484_));
 XOR2_X2 _30650_ (.A(_05369_),
    .B(_05484_),
    .Z(_05485_));
 NOR2_X2 _30651_ (.A1(_16726_),
    .A2(_16725_),
    .ZN(_05486_));
 NOR2_X1 _30652_ (.A1(_16724_),
    .A2(_16723_),
    .ZN(_05487_));
 CLKBUF_X2 _30653_ (.A(_05487_),
    .Z(_05488_));
 AND2_X2 _30654_ (.A1(_05486_),
    .A2(_05488_),
    .ZN(_05490_));
 CLKBUF_X2 _30655_ (.A(_05490_),
    .Z(_05491_));
 AND2_X1 _30656_ (.A1(_16721_),
    .A2(_16722_),
    .ZN(_05492_));
 CLKBUF_X2 _30657_ (.A(_05492_),
    .Z(_05493_));
 INV_X2 _30658_ (.A(_16720_),
    .ZN(_05494_));
 NOR2_X2 _30659_ (.A1(_05494_),
    .A2(_16719_),
    .ZN(_05495_));
 CLKBUF_X2 _30660_ (.A(_05495_),
    .Z(_05496_));
 INV_X1 _30661_ (.A(_16719_),
    .ZN(_05497_));
 NOR2_X2 _30662_ (.A1(_05497_),
    .A2(_16720_),
    .ZN(_05498_));
 BUF_X2 _30663_ (.A(_05498_),
    .Z(_05499_));
 OAI211_X1 _30664_ (.A(_05491_),
    .B(_05493_),
    .C1(_05496_),
    .C2(_05499_),
    .ZN(_05501_));
 INV_X1 _30665_ (.A(_16722_),
    .ZN(_05502_));
 NOR2_X1 _30666_ (.A1(_05502_),
    .A2(_16721_),
    .ZN(_05503_));
 CLKBUF_X2 _30667_ (.A(_05503_),
    .Z(_05504_));
 CLKBUF_X2 _30668_ (.A(_05504_),
    .Z(_05505_));
 CLKBUF_X2 _30669_ (.A(_05486_),
    .Z(_05506_));
 NAND4_X1 _30670_ (.A1(_05505_),
    .A2(_05499_),
    .A3(_05506_),
    .A4(_05488_),
    .ZN(_05507_));
 AND2_X2 _30671_ (.A1(_05503_),
    .A2(_16720_),
    .ZN(_05508_));
 INV_X2 _30672_ (.A(_05508_),
    .ZN(_05509_));
 INV_X1 _30673_ (.A(_05490_),
    .ZN(_05510_));
 OAI211_X1 _30674_ (.A(_05501_),
    .B(_05507_),
    .C1(_05509_),
    .C2(_05510_),
    .ZN(_05512_));
 NOR2_X1 _30675_ (.A1(_16721_),
    .A2(_16722_),
    .ZN(_05513_));
 CLKBUF_X2 _30676_ (.A(_05513_),
    .Z(_05514_));
 CLKBUF_X2 _30677_ (.A(_16720_),
    .Z(_05515_));
 AND2_X1 _30678_ (.A1(_05514_),
    .A2(_05515_),
    .ZN(_05516_));
 AND2_X1 _30679_ (.A1(_05491_),
    .A2(_05516_),
    .ZN(_05517_));
 INV_X1 _30680_ (.A(_16721_),
    .ZN(_05518_));
 NOR2_X1 _30681_ (.A1(_05518_),
    .A2(_16722_),
    .ZN(_05519_));
 AND2_X1 _30682_ (.A1(_05519_),
    .A2(_05515_),
    .ZN(_05520_));
 CLKBUF_X2 _30683_ (.A(_05520_),
    .Z(_05521_));
 AND2_X1 _30684_ (.A1(_05521_),
    .A2(_05491_),
    .ZN(_05523_));
 CLKBUF_X2 _30685_ (.A(_05519_),
    .Z(_05524_));
 CLKBUF_X2 _30686_ (.A(_05524_),
    .Z(_05525_));
 AND3_X1 _30687_ (.A1(_05491_),
    .A2(_05525_),
    .A3(_05499_),
    .ZN(_05526_));
 NOR4_X1 _30688_ (.A1(_05512_),
    .A2(_05517_),
    .A3(_05523_),
    .A4(_05526_),
    .ZN(_05527_));
 INV_X1 _30689_ (.A(_16724_),
    .ZN(_05528_));
 AND2_X1 _30690_ (.A1(_05528_),
    .A2(_16723_),
    .ZN(_05529_));
 AND2_X1 _30691_ (.A1(_05529_),
    .A2(_05486_),
    .ZN(_05530_));
 NOR2_X2 _30692_ (.A1(_16720_),
    .A2(_16719_),
    .ZN(_05531_));
 INV_X2 _30693_ (.A(_05531_),
    .ZN(_05532_));
 AND2_X1 _30694_ (.A1(_05532_),
    .A2(_05519_),
    .ZN(_05534_));
 AND2_X2 _30695_ (.A1(_16720_),
    .A2(_16719_),
    .ZN(_05535_));
 INV_X1 _30696_ (.A(_05535_),
    .ZN(_05536_));
 CLKBUF_X2 _30697_ (.A(_05536_),
    .Z(_05537_));
 AND3_X1 _30698_ (.A1(_05530_),
    .A2(_05534_),
    .A3(_05537_),
    .ZN(_05538_));
 OAI21_X1 _30699_ (.A(_05504_),
    .B1(_05494_),
    .B2(_16719_),
    .ZN(_05539_));
 NOR2_X1 _30700_ (.A1(_05539_),
    .A2(_05499_),
    .ZN(_05540_));
 BUF_X2 _30701_ (.A(_05530_),
    .Z(_05541_));
 AND2_X1 _30702_ (.A1(_05540_),
    .A2(_05541_),
    .ZN(_05542_));
 BUF_X2 _30703_ (.A(_05516_),
    .Z(_05543_));
 AOI211_X1 _30704_ (.A(_05538_),
    .B(_05542_),
    .C1(_05541_),
    .C2(_05543_),
    .ZN(_05545_));
 NOR2_X1 _30705_ (.A1(_05528_),
    .A2(_16723_),
    .ZN(_05546_));
 AND2_X1 _30706_ (.A1(_05546_),
    .A2(_05486_),
    .ZN(_05547_));
 INV_X1 _30707_ (.A(_05547_),
    .ZN(_05548_));
 NAND2_X1 _30708_ (.A1(_05536_),
    .A2(_05514_),
    .ZN(_05549_));
 NOR2_X1 _30709_ (.A1(_05548_),
    .A2(_05549_),
    .ZN(_05550_));
 INV_X1 _30710_ (.A(_05550_),
    .ZN(_05551_));
 AND3_X1 _30711_ (.A1(_05547_),
    .A2(_05504_),
    .A3(_05532_),
    .ZN(_05552_));
 INV_X1 _30712_ (.A(_05552_),
    .ZN(_05553_));
 BUF_X2 _30713_ (.A(_05547_),
    .Z(_05554_));
 NAND3_X1 _30714_ (.A1(_05534_),
    .A2(_05554_),
    .A3(_05537_),
    .ZN(_05556_));
 AND2_X2 _30715_ (.A1(_05493_),
    .A2(_05531_),
    .ZN(_05557_));
 AND2_X1 _30716_ (.A1(_05493_),
    .A2(_05515_),
    .ZN(_05558_));
 OAI21_X1 _30717_ (.A(_05554_),
    .B1(_05557_),
    .B2(_05558_),
    .ZN(_05559_));
 AND4_X1 _30718_ (.A1(_05551_),
    .A2(_05553_),
    .A3(_05556_),
    .A4(_05559_),
    .ZN(_05560_));
 AND2_X1 _30719_ (.A1(_16724_),
    .A2(_16723_),
    .ZN(_05561_));
 AND2_X1 _30720_ (.A1(_05561_),
    .A2(_05486_),
    .ZN(_05562_));
 INV_X1 _30721_ (.A(_05562_),
    .ZN(_05563_));
 AND2_X2 _30722_ (.A1(_05496_),
    .A2(_05519_),
    .ZN(_05564_));
 INV_X1 _30723_ (.A(_05564_),
    .ZN(_05565_));
 CLKBUF_X2 _30724_ (.A(_05514_),
    .Z(_05567_));
 NAND2_X1 _30725_ (.A1(_05532_),
    .A2(_05567_),
    .ZN(_05568_));
 AOI21_X1 _30726_ (.A(_05563_),
    .B1(_05565_),
    .B2(_05568_),
    .ZN(_05569_));
 AND2_X2 _30727_ (.A1(_05492_),
    .A2(_05535_),
    .ZN(_05570_));
 AND2_X1 _30728_ (.A1(_05570_),
    .A2(_05562_),
    .ZN(_05571_));
 CLKBUF_X2 _30729_ (.A(_05531_),
    .Z(_05572_));
 AND3_X1 _30730_ (.A1(_05562_),
    .A2(_05505_),
    .A3(_05572_),
    .ZN(_05573_));
 NAND2_X1 _30731_ (.A1(_05494_),
    .A2(_16722_),
    .ZN(_05574_));
 NOR2_X2 _30732_ (.A1(_05574_),
    .A2(_05518_),
    .ZN(_05575_));
 AND2_X1 _30733_ (.A1(_05562_),
    .A2(_05575_),
    .ZN(_05576_));
 NOR4_X1 _30734_ (.A1(_05569_),
    .A2(_05571_),
    .A3(_05573_),
    .A4(_05576_),
    .ZN(_05578_));
 AND4_X1 _30735_ (.A1(_05527_),
    .A2(_05545_),
    .A3(_05560_),
    .A4(_05578_),
    .ZN(_05579_));
 INV_X1 _30736_ (.A(_16725_),
    .ZN(_05580_));
 NOR2_X1 _30737_ (.A1(_05580_),
    .A2(_16726_),
    .ZN(_05581_));
 AND2_X1 _30738_ (.A1(_05581_),
    .A2(_05488_),
    .ZN(_05582_));
 BUF_X2 _30739_ (.A(_05582_),
    .Z(_05583_));
 AND2_X1 _30740_ (.A1(_05514_),
    .A2(_05494_),
    .ZN(_05584_));
 INV_X1 _30741_ (.A(_05584_),
    .ZN(_05585_));
 INV_X1 _30742_ (.A(_05525_),
    .ZN(_05586_));
 OAI21_X1 _30743_ (.A(_05585_),
    .B1(_05586_),
    .B2(_05532_),
    .ZN(_05587_));
 CLKBUF_X2 _30744_ (.A(_05493_),
    .Z(_05589_));
 CLKBUF_X2 _30745_ (.A(_05497_),
    .Z(_05590_));
 OAI21_X1 _30746_ (.A(_05589_),
    .B1(_05494_),
    .B2(_05590_),
    .ZN(_05591_));
 INV_X1 _30747_ (.A(_05505_),
    .ZN(_05592_));
 CLKBUF_X2 _30748_ (.A(_05590_),
    .Z(_05593_));
 OAI21_X1 _30749_ (.A(_05591_),
    .B1(_05592_),
    .B2(_05593_),
    .ZN(_05594_));
 OAI21_X1 _30750_ (.A(_05583_),
    .B1(_05587_),
    .B2(_05594_),
    .ZN(_05595_));
 CLKBUF_X2 _30751_ (.A(_05546_),
    .Z(_05596_));
 AND2_X1 _30752_ (.A1(_05596_),
    .A2(_05581_),
    .ZN(_05597_));
 INV_X1 _30753_ (.A(_05597_),
    .ZN(_05598_));
 NOR2_X1 _30754_ (.A1(_05598_),
    .A2(_05539_),
    .ZN(_05600_));
 AND2_X1 _30755_ (.A1(_05514_),
    .A2(_16719_),
    .ZN(_05601_));
 INV_X1 _30756_ (.A(_05601_),
    .ZN(_05602_));
 AOI21_X1 _30757_ (.A(_05598_),
    .B1(_05586_),
    .B2(_05602_),
    .ZN(_05603_));
 AND2_X1 _30758_ (.A1(_05495_),
    .A2(_05492_),
    .ZN(_05604_));
 BUF_X2 _30759_ (.A(_05604_),
    .Z(_05605_));
 CLKBUF_X2 _30760_ (.A(_05597_),
    .Z(_05606_));
 AOI211_X1 _30761_ (.A(_05600_),
    .B(_05603_),
    .C1(_05605_),
    .C2(_05606_),
    .ZN(_05607_));
 AND2_X1 _30762_ (.A1(_05529_),
    .A2(_05581_),
    .ZN(_05608_));
 BUF_X2 _30763_ (.A(_05608_),
    .Z(_05609_));
 CLKBUF_X2 _30764_ (.A(_16719_),
    .Z(_05611_));
 AND2_X1 _30765_ (.A1(_05505_),
    .A2(_05611_),
    .ZN(_05612_));
 OAI21_X1 _30766_ (.A(_05609_),
    .B1(_05612_),
    .B2(_05570_),
    .ZN(_05613_));
 AND2_X1 _30767_ (.A1(_05609_),
    .A2(_05521_),
    .ZN(_05614_));
 INV_X1 _30768_ (.A(_05614_),
    .ZN(_05615_));
 BUF_X2 _30769_ (.A(_05584_),
    .Z(_05616_));
 NAND2_X1 _30770_ (.A1(_05609_),
    .A2(_05616_),
    .ZN(_05617_));
 AND2_X1 _30771_ (.A1(_05535_),
    .A2(_05514_),
    .ZN(_05618_));
 BUF_X2 _30772_ (.A(_05618_),
    .Z(_05619_));
 NAND2_X1 _30773_ (.A1(_05609_),
    .A2(_05619_),
    .ZN(_05620_));
 AND4_X1 _30774_ (.A1(_05613_),
    .A2(_05615_),
    .A3(_05617_),
    .A4(_05620_),
    .ZN(_05622_));
 NOR2_X1 _30775_ (.A1(_05497_),
    .A2(_16722_),
    .ZN(_05623_));
 AND2_X1 _30776_ (.A1(_05623_),
    .A2(_16721_),
    .ZN(_05624_));
 AND2_X1 _30777_ (.A1(_05581_),
    .A2(_05561_),
    .ZN(_05625_));
 BUF_X2 _30778_ (.A(_05625_),
    .Z(_05626_));
 NAND2_X1 _30779_ (.A1(_05624_),
    .A2(_05626_),
    .ZN(_05627_));
 AND2_X1 _30780_ (.A1(_05498_),
    .A2(_05493_),
    .ZN(_05628_));
 OAI21_X1 _30781_ (.A(_05625_),
    .B1(_05605_),
    .B2(_05628_),
    .ZN(_05629_));
 OAI21_X1 _30782_ (.A(_05625_),
    .B1(_05618_),
    .B2(_05616_),
    .ZN(_05630_));
 AND2_X1 _30783_ (.A1(_05504_),
    .A2(_05535_),
    .ZN(_05631_));
 BUF_X2 _30784_ (.A(_05631_),
    .Z(_05633_));
 NAND2_X1 _30785_ (.A1(_05625_),
    .A2(_05633_),
    .ZN(_05634_));
 AND4_X1 _30786_ (.A1(_05627_),
    .A2(_05629_),
    .A3(_05630_),
    .A4(_05634_),
    .ZN(_05635_));
 AND4_X1 _30787_ (.A1(_05595_),
    .A2(_05607_),
    .A3(_05622_),
    .A4(_05635_),
    .ZN(_05636_));
 AND2_X1 _30788_ (.A1(_05580_),
    .A2(_16726_),
    .ZN(_05637_));
 CLKBUF_X2 _30789_ (.A(_05637_),
    .Z(_05638_));
 OAI211_X1 _30790_ (.A(_05596_),
    .B(_05638_),
    .C1(_05570_),
    .C2(_05575_),
    .ZN(_05639_));
 NAND4_X1 _30791_ (.A1(_05638_),
    .A2(_05505_),
    .A3(_05499_),
    .A4(_05596_),
    .ZN(_05640_));
 AND2_X1 _30792_ (.A1(_05639_),
    .A2(_05640_),
    .ZN(_05641_));
 AND2_X2 _30793_ (.A1(_05637_),
    .A2(_05529_),
    .ZN(_05642_));
 AND2_X2 _30794_ (.A1(_05496_),
    .A2(_05514_),
    .ZN(_05644_));
 AND2_X1 _30795_ (.A1(_05498_),
    .A2(_05514_),
    .ZN(_05645_));
 CLKBUF_X2 _30796_ (.A(_05645_),
    .Z(_05646_));
 OAI21_X1 _30797_ (.A(_05642_),
    .B1(_05644_),
    .B2(_05646_),
    .ZN(_05647_));
 INV_X1 _30798_ (.A(_05558_),
    .ZN(_05648_));
 INV_X2 _30799_ (.A(_05642_),
    .ZN(_05649_));
 OAI21_X1 _30800_ (.A(_05647_),
    .B1(_05648_),
    .B2(_05649_),
    .ZN(_05650_));
 AND2_X2 _30801_ (.A1(_05637_),
    .A2(_05487_),
    .ZN(_05651_));
 INV_X1 _30802_ (.A(_05651_),
    .ZN(_05652_));
 INV_X1 _30803_ (.A(_05612_),
    .ZN(_05653_));
 NAND2_X1 _30804_ (.A1(_05532_),
    .A2(_05493_),
    .ZN(_05655_));
 AOI21_X1 _30805_ (.A(_05652_),
    .B1(_05653_),
    .B2(_05655_),
    .ZN(_05656_));
 INV_X1 _30806_ (.A(_05495_),
    .ZN(_05657_));
 NAND2_X1 _30807_ (.A1(_05657_),
    .A2(_05524_),
    .ZN(_05658_));
 NOR2_X1 _30808_ (.A1(_05652_),
    .A2(_05658_),
    .ZN(_05659_));
 AND4_X1 _30809_ (.A1(_05590_),
    .A2(_05638_),
    .A3(_05567_),
    .A4(_05488_),
    .ZN(_05660_));
 NOR4_X1 _30810_ (.A1(_05650_),
    .A2(_05656_),
    .A3(_05659_),
    .A4(_05660_),
    .ZN(_05661_));
 AND2_X1 _30811_ (.A1(_05637_),
    .A2(_05561_),
    .ZN(_05662_));
 INV_X1 _30812_ (.A(_05662_),
    .ZN(_05663_));
 INV_X1 _30813_ (.A(_05498_),
    .ZN(_05664_));
 CLKBUF_X2 _30814_ (.A(_05664_),
    .Z(_05666_));
 NAND2_X1 _30815_ (.A1(_05666_),
    .A2(_05567_),
    .ZN(_05667_));
 NOR2_X1 _30816_ (.A1(_05663_),
    .A2(_05667_),
    .ZN(_05668_));
 NOR2_X1 _30817_ (.A1(_05663_),
    .A2(_05658_),
    .ZN(_05669_));
 BUF_X2 _30818_ (.A(_05662_),
    .Z(_05670_));
 AOI211_X1 _30819_ (.A(_05668_),
    .B(_05669_),
    .C1(_05557_),
    .C2(_05670_),
    .ZN(_05671_));
 AND2_X1 _30820_ (.A1(_05637_),
    .A2(_05596_),
    .ZN(_05672_));
 BUF_X2 _30821_ (.A(_05672_),
    .Z(_05673_));
 AND2_X1 _30822_ (.A1(_05524_),
    .A2(_05531_),
    .ZN(_05674_));
 AND2_X1 _30823_ (.A1(_05673_),
    .A2(_05674_),
    .ZN(_05675_));
 INV_X1 _30824_ (.A(_05675_),
    .ZN(_05677_));
 AND4_X1 _30825_ (.A1(_05641_),
    .A2(_05661_),
    .A3(_05671_),
    .A4(_05677_),
    .ZN(_05678_));
 AND2_X2 _30826_ (.A1(_16726_),
    .A2(_16725_),
    .ZN(_05679_));
 AND2_X1 _30827_ (.A1(_05546_),
    .A2(_05679_),
    .ZN(_05680_));
 CLKBUF_X2 _30828_ (.A(_05680_),
    .Z(_05681_));
 INV_X1 _30829_ (.A(_05681_),
    .ZN(_05682_));
 OAI21_X1 _30830_ (.A(_05504_),
    .B1(_05515_),
    .B2(_05590_),
    .ZN(_05683_));
 NOR2_X1 _30831_ (.A1(_05682_),
    .A2(_05683_),
    .ZN(_05684_));
 INV_X1 _30832_ (.A(_05513_),
    .ZN(_05685_));
 NOR2_X1 _30833_ (.A1(_05685_),
    .A2(_05495_),
    .ZN(_05686_));
 AND3_X1 _30834_ (.A1(_05681_),
    .A2(_05686_),
    .A3(_05664_),
    .ZN(_05688_));
 AND2_X1 _30835_ (.A1(_05519_),
    .A2(_05494_),
    .ZN(_05689_));
 CLKBUF_X2 _30836_ (.A(_05689_),
    .Z(_05690_));
 AND2_X1 _30837_ (.A1(_05690_),
    .A2(_05681_),
    .ZN(_05691_));
 AND2_X1 _30838_ (.A1(_05493_),
    .A2(_16719_),
    .ZN(_05692_));
 AND3_X1 _30839_ (.A1(_05692_),
    .A2(_05679_),
    .A3(_05596_),
    .ZN(_05693_));
 OR4_X1 _30840_ (.A1(_05684_),
    .A2(_05688_),
    .A3(_05691_),
    .A4(_05693_),
    .ZN(_05694_));
 AND2_X1 _30841_ (.A1(_05529_),
    .A2(_05679_),
    .ZN(_05695_));
 BUF_X2 _30842_ (.A(_05695_),
    .Z(_05696_));
 AND2_X1 _30843_ (.A1(_05519_),
    .A2(_05498_),
    .ZN(_05697_));
 BUF_X2 _30844_ (.A(_05697_),
    .Z(_05699_));
 OAI21_X1 _30845_ (.A(_05696_),
    .B1(_05699_),
    .B2(_05644_),
    .ZN(_05700_));
 BUF_X2 _30846_ (.A(_05628_),
    .Z(_05701_));
 OAI21_X1 _30847_ (.A(_05696_),
    .B1(_05605_),
    .B2(_05701_),
    .ZN(_05702_));
 BUF_X2 _30848_ (.A(_05508_),
    .Z(_05703_));
 NOR2_X2 _30849_ (.A1(_05574_),
    .A2(_16721_),
    .ZN(_05704_));
 BUF_X2 _30850_ (.A(_05704_),
    .Z(_05705_));
 OAI21_X1 _30851_ (.A(_05696_),
    .B1(_05703_),
    .B2(_05705_),
    .ZN(_05706_));
 NAND3_X1 _30852_ (.A1(_05700_),
    .A2(_05702_),
    .A3(_05706_),
    .ZN(_05707_));
 AND2_X1 _30853_ (.A1(_05679_),
    .A2(_05487_),
    .ZN(_05708_));
 BUF_X2 _30854_ (.A(_05708_),
    .Z(_05710_));
 BUF_X2 _30855_ (.A(_05494_),
    .Z(_05711_));
 OAI211_X1 _30856_ (.A(_05710_),
    .B(_05589_),
    .C1(_05711_),
    .C2(_05593_),
    .ZN(_05712_));
 BUF_X2 _30857_ (.A(_05496_),
    .Z(_05713_));
 CLKBUF_X2 _30858_ (.A(_05679_),
    .Z(_05714_));
 CLKBUF_X2 _30859_ (.A(_05567_),
    .Z(_05715_));
 CLKBUF_X2 _30860_ (.A(_05488_),
    .Z(_05716_));
 NAND4_X1 _30861_ (.A1(_05713_),
    .A2(_05714_),
    .A3(_05715_),
    .A4(_05716_),
    .ZN(_05717_));
 INV_X1 _30862_ (.A(_05710_),
    .ZN(_05718_));
 OAI211_X1 _30863_ (.A(_05712_),
    .B(_05717_),
    .C1(_05718_),
    .C2(_05653_),
    .ZN(_05719_));
 AND2_X2 _30864_ (.A1(_05679_),
    .A2(_05561_),
    .ZN(_05721_));
 BUF_X2 _30865_ (.A(_05721_),
    .Z(_05722_));
 OAI21_X1 _30866_ (.A(_05722_),
    .B1(_05508_),
    .B2(_05705_),
    .ZN(_05723_));
 OAI211_X1 _30867_ (.A(_05721_),
    .B(_05715_),
    .C1(_05515_),
    .C2(_05611_),
    .ZN(_05724_));
 NAND2_X1 _30868_ (.A1(_05674_),
    .A2(_05722_),
    .ZN(_05725_));
 NAND3_X1 _30869_ (.A1(_05721_),
    .A2(_05589_),
    .A3(_05713_),
    .ZN(_05726_));
 NAND4_X1 _30870_ (.A1(_05723_),
    .A2(_05724_),
    .A3(_05725_),
    .A4(_05726_),
    .ZN(_05727_));
 NOR4_X1 _30871_ (.A1(_05694_),
    .A2(_05707_),
    .A3(_05719_),
    .A4(_05727_),
    .ZN(_05728_));
 NAND4_X1 _30872_ (.A1(_05579_),
    .A2(_05636_),
    .A3(_05678_),
    .A4(_05728_),
    .ZN(_05729_));
 OAI21_X1 _30873_ (.A(_05502_),
    .B1(_05532_),
    .B2(_16721_),
    .ZN(_05730_));
 AND3_X1 _30874_ (.A1(_05506_),
    .A2(_05488_),
    .A3(_05502_),
    .ZN(_05732_));
 AND2_X1 _30875_ (.A1(_05730_),
    .A2(_05732_),
    .ZN(_05733_));
 OR2_X2 _30876_ (.A1(_05729_),
    .A2(_05733_),
    .ZN(_05734_));
 XNOR2_X1 _30877_ (.A(_05734_),
    .B(_14166_),
    .ZN(_05735_));
 XNOR2_X1 _30878_ (.A(_05485_),
    .B(_05735_),
    .ZN(_05736_));
 INV_X1 _30879_ (.A(_16801_),
    .ZN(_05737_));
 NOR2_X1 _30880_ (.A1(_05737_),
    .A2(_16802_),
    .ZN(_05738_));
 CLKBUF_X2 _30881_ (.A(_05738_),
    .Z(_05739_));
 INV_X1 _30882_ (.A(_05739_),
    .ZN(_05740_));
 INV_X1 _30883_ (.A(_16800_),
    .ZN(_05741_));
 NOR2_X2 _30884_ (.A1(_05741_),
    .A2(_16799_),
    .ZN(_05743_));
 NOR2_X2 _30885_ (.A1(_05740_),
    .A2(_05743_),
    .ZN(_05744_));
 INV_X1 _30886_ (.A(_16799_),
    .ZN(_05745_));
 NOR2_X2 _30887_ (.A1(_05745_),
    .A2(_16800_),
    .ZN(_05746_));
 INV_X1 _30888_ (.A(_05746_),
    .ZN(_05747_));
 NOR2_X2 _30889_ (.A1(_16804_),
    .A2(_16803_),
    .ZN(_05748_));
 NOR2_X2 _30890_ (.A1(_16805_),
    .A2(_16806_),
    .ZN(_05749_));
 AND2_X1 _30891_ (.A1(_05748_),
    .A2(_05749_),
    .ZN(_05750_));
 BUF_X2 _30892_ (.A(_05750_),
    .Z(_05751_));
 NAND3_X1 _30893_ (.A1(_05744_),
    .A2(_05747_),
    .A3(_05751_),
    .ZN(_05752_));
 INV_X1 _30894_ (.A(_16804_),
    .ZN(_05754_));
 AND2_X1 _30895_ (.A1(_05754_),
    .A2(_16803_),
    .ZN(_05755_));
 CLKBUF_X2 _30896_ (.A(_05755_),
    .Z(_05756_));
 AND2_X1 _30897_ (.A1(_05756_),
    .A2(_05749_),
    .ZN(_05757_));
 NOR2_X1 _30898_ (.A1(_16802_),
    .A2(_16801_),
    .ZN(_05758_));
 CLKBUF_X2 _30899_ (.A(_05758_),
    .Z(_05759_));
 AND2_X1 _30900_ (.A1(_05759_),
    .A2(_05741_),
    .ZN(_05760_));
 AND2_X1 _30901_ (.A1(_05757_),
    .A2(_05760_),
    .ZN(_05761_));
 NOR2_X1 _30902_ (.A1(_16799_),
    .A2(_16800_),
    .ZN(_05762_));
 CLKBUF_X2 _30903_ (.A(_05762_),
    .Z(_05763_));
 AND2_X1 _30904_ (.A1(_05738_),
    .A2(_05763_),
    .ZN(_05765_));
 INV_X1 _30905_ (.A(_05765_),
    .ZN(_05766_));
 AND2_X2 _30906_ (.A1(_16799_),
    .A2(_16800_),
    .ZN(_05767_));
 AND2_X1 _30907_ (.A1(_05738_),
    .A2(_05767_),
    .ZN(_05768_));
 INV_X1 _30908_ (.A(_05768_),
    .ZN(_05769_));
 NAND2_X1 _30909_ (.A1(_05766_),
    .A2(_05769_),
    .ZN(_05770_));
 CLKBUF_X2 _30910_ (.A(_05757_),
    .Z(_05771_));
 AND2_X1 _30911_ (.A1(_05770_),
    .A2(_05771_),
    .ZN(_05772_));
 AND2_X1 _30912_ (.A1(_05743_),
    .A2(_05758_),
    .ZN(_05773_));
 BUF_X2 _30913_ (.A(_05757_),
    .Z(_05774_));
 AOI211_X1 _30914_ (.A(_05761_),
    .B(_05772_),
    .C1(_05773_),
    .C2(_05774_),
    .ZN(_05776_));
 AND2_X1 _30915_ (.A1(_16802_),
    .A2(_16801_),
    .ZN(_05777_));
 CLKBUF_X2 _30916_ (.A(_05777_),
    .Z(_05778_));
 CLKBUF_X2 _30917_ (.A(_05778_),
    .Z(_05779_));
 BUF_X2 _30918_ (.A(_05745_),
    .Z(_05780_));
 BUF_X2 _30919_ (.A(_05741_),
    .Z(_05781_));
 OAI211_X1 _30920_ (.A(_05751_),
    .B(_05779_),
    .C1(_05780_),
    .C2(_05781_),
    .ZN(_05782_));
 AND2_X2 _30921_ (.A1(_05777_),
    .A2(_05767_),
    .ZN(_05783_));
 NAND2_X1 _30922_ (.A1(_05757_),
    .A2(_05783_),
    .ZN(_05784_));
 INV_X1 _30923_ (.A(_16802_),
    .ZN(_05785_));
 NOR2_X1 _30924_ (.A1(_05785_),
    .A2(_16801_),
    .ZN(_05787_));
 AND2_X1 _30925_ (.A1(_05787_),
    .A2(_05741_),
    .ZN(_05788_));
 CLKBUF_X2 _30926_ (.A(_05788_),
    .Z(_05789_));
 NAND2_X1 _30927_ (.A1(_05771_),
    .A2(_05789_),
    .ZN(_05790_));
 NOR2_X1 _30928_ (.A1(_05741_),
    .A2(_16801_),
    .ZN(_05791_));
 AND2_X1 _30929_ (.A1(_05791_),
    .A2(_16802_),
    .ZN(_05792_));
 NAND2_X1 _30930_ (.A1(_05757_),
    .A2(_05792_),
    .ZN(_05793_));
 AND2_X1 _30931_ (.A1(_05778_),
    .A2(_05741_),
    .ZN(_05794_));
 NAND2_X1 _30932_ (.A1(_05771_),
    .A2(_05794_),
    .ZN(_05795_));
 AND4_X1 _30933_ (.A1(_05784_),
    .A2(_05790_),
    .A3(_05793_),
    .A4(_05795_),
    .ZN(_05796_));
 AND4_X1 _30934_ (.A1(_05752_),
    .A2(_05776_),
    .A3(_05782_),
    .A4(_05796_),
    .ZN(_05798_));
 INV_X1 _30935_ (.A(_16805_),
    .ZN(_05799_));
 NOR2_X1 _30936_ (.A1(_05799_),
    .A2(_16806_),
    .ZN(_05800_));
 AND2_X1 _30937_ (.A1(_16804_),
    .A2(_16803_),
    .ZN(_05801_));
 CLKBUF_X2 _30938_ (.A(_05801_),
    .Z(_05802_));
 AND2_X1 _30939_ (.A1(_05800_),
    .A2(_05802_),
    .ZN(_05803_));
 AND2_X1 _30940_ (.A1(_05759_),
    .A2(_16799_),
    .ZN(_05804_));
 AND2_X1 _30941_ (.A1(_05803_),
    .A2(_05804_),
    .ZN(_05805_));
 INV_X1 _30942_ (.A(_05805_),
    .ZN(_05806_));
 BUF_X2 _30943_ (.A(_05768_),
    .Z(_05807_));
 CLKBUF_X2 _30944_ (.A(_05803_),
    .Z(_05809_));
 NAND2_X1 _30945_ (.A1(_05807_),
    .A2(_05809_),
    .ZN(_05810_));
 AND2_X1 _30946_ (.A1(_05738_),
    .A2(_05741_),
    .ZN(_05811_));
 INV_X1 _30947_ (.A(_05811_),
    .ZN(_05812_));
 INV_X1 _30948_ (.A(_05809_),
    .ZN(_05813_));
 OAI211_X1 _30949_ (.A(_05806_),
    .B(_05810_),
    .C1(_05812_),
    .C2(_05813_),
    .ZN(_05814_));
 AND2_X1 _30950_ (.A1(_05809_),
    .A2(_05789_),
    .ZN(_05815_));
 AND2_X1 _30951_ (.A1(_05787_),
    .A2(_05743_),
    .ZN(_05816_));
 BUF_X2 _30952_ (.A(_05816_),
    .Z(_05817_));
 AND2_X1 _30953_ (.A1(_05817_),
    .A2(_05803_),
    .ZN(_05818_));
 OR2_X1 _30954_ (.A1(_05815_),
    .A2(_05818_),
    .ZN(_05820_));
 INV_X1 _30955_ (.A(_05762_),
    .ZN(_05821_));
 NAND2_X1 _30956_ (.A1(_05821_),
    .A2(_05777_),
    .ZN(_05822_));
 INV_X1 _30957_ (.A(_05822_),
    .ZN(_05823_));
 AND2_X1 _30958_ (.A1(_05823_),
    .A2(_05803_),
    .ZN(_05824_));
 NOR2_X2 _30959_ (.A1(_05754_),
    .A2(_16803_),
    .ZN(_05825_));
 AND2_X1 _30960_ (.A1(_05800_),
    .A2(_05825_),
    .ZN(_05826_));
 BUF_X2 _30961_ (.A(_05826_),
    .Z(_05827_));
 BUF_X2 _30962_ (.A(_05827_),
    .Z(_05828_));
 CLKBUF_X2 _30963_ (.A(_05760_),
    .Z(_05829_));
 AND2_X2 _30964_ (.A1(_05758_),
    .A2(_16800_),
    .ZN(_05831_));
 OAI21_X1 _30965_ (.A(_05828_),
    .B1(_05829_),
    .B2(_05831_),
    .ZN(_05832_));
 CLKBUF_X2 _30966_ (.A(_05787_),
    .Z(_05833_));
 AND2_X2 _30967_ (.A1(_05833_),
    .A2(_05746_),
    .ZN(_05834_));
 NAND2_X1 _30968_ (.A1(_05834_),
    .A2(_05827_),
    .ZN(_05835_));
 NAND2_X1 _30969_ (.A1(_05827_),
    .A2(_05807_),
    .ZN(_05836_));
 AND2_X1 _30970_ (.A1(_05777_),
    .A2(_16800_),
    .ZN(_05837_));
 NAND2_X1 _30971_ (.A1(_05827_),
    .A2(_05837_),
    .ZN(_05838_));
 NAND4_X1 _30972_ (.A1(_05832_),
    .A2(_05835_),
    .A3(_05836_),
    .A4(_05838_),
    .ZN(_05839_));
 NOR4_X1 _30973_ (.A1(_05814_),
    .A2(_05820_),
    .A3(_05824_),
    .A4(_05839_),
    .ZN(_05840_));
 AND2_X1 _30974_ (.A1(_05756_),
    .A2(_05800_),
    .ZN(_05842_));
 BUF_X2 _30975_ (.A(_05842_),
    .Z(_05843_));
 NOR3_X1 _30976_ (.A1(_05762_),
    .A2(_05785_),
    .A3(_16801_),
    .ZN(_05844_));
 INV_X1 _30977_ (.A(_05767_),
    .ZN(_05845_));
 AND2_X1 _30978_ (.A1(_05844_),
    .A2(_05845_),
    .ZN(_05846_));
 OAI21_X1 _30979_ (.A(_05843_),
    .B1(_05846_),
    .B2(_05783_),
    .ZN(_05847_));
 BUF_X2 _30980_ (.A(_05756_),
    .Z(_05848_));
 CLKBUF_X2 _30981_ (.A(_05800_),
    .Z(_05849_));
 BUF_X2 _30982_ (.A(_16799_),
    .Z(_05850_));
 BUF_X2 _30983_ (.A(_05759_),
    .Z(_05851_));
 NAND4_X1 _30984_ (.A1(_05848_),
    .A2(_05849_),
    .A3(_05850_),
    .A4(_05851_),
    .ZN(_05853_));
 AND2_X1 _30985_ (.A1(_05746_),
    .A2(_05738_),
    .ZN(_05854_));
 BUF_X2 _30986_ (.A(_05854_),
    .Z(_05855_));
 AND2_X1 _30987_ (.A1(_05743_),
    .A2(_05738_),
    .ZN(_05856_));
 BUF_X2 _30988_ (.A(_05856_),
    .Z(_05857_));
 OAI21_X1 _30989_ (.A(_05843_),
    .B1(_05855_),
    .B2(_05857_),
    .ZN(_05858_));
 AND3_X1 _30990_ (.A1(_05847_),
    .A2(_05853_),
    .A3(_05858_),
    .ZN(_05859_));
 AND2_X1 _30991_ (.A1(_05849_),
    .A2(_05748_),
    .ZN(_05860_));
 BUF_X2 _30992_ (.A(_05860_),
    .Z(_05861_));
 AND2_X1 _30993_ (.A1(_05746_),
    .A2(_05759_),
    .ZN(_05862_));
 CLKBUF_X2 _30994_ (.A(_05862_),
    .Z(_05864_));
 OAI21_X1 _30995_ (.A(_05861_),
    .B1(_05807_),
    .B2(_05864_),
    .ZN(_05865_));
 CLKBUF_X2 _30996_ (.A(_05792_),
    .Z(_05866_));
 AND2_X2 _30997_ (.A1(_05778_),
    .A2(_16799_),
    .ZN(_05867_));
 OAI21_X1 _30998_ (.A(_05861_),
    .B1(_05866_),
    .B2(_05867_),
    .ZN(_05868_));
 AND3_X1 _30999_ (.A1(_05859_),
    .A2(_05865_),
    .A3(_05868_),
    .ZN(_05869_));
 AND2_X1 _31000_ (.A1(_05825_),
    .A2(_05749_),
    .ZN(_05870_));
 INV_X1 _31001_ (.A(_05870_),
    .ZN(_05871_));
 CLKBUF_X2 _31002_ (.A(_05845_),
    .Z(_05872_));
 NAND2_X1 _31003_ (.A1(_05872_),
    .A2(_05759_),
    .ZN(_05873_));
 NOR2_X1 _31004_ (.A1(_05871_),
    .A2(_05873_),
    .ZN(_05875_));
 AND2_X1 _31005_ (.A1(_05739_),
    .A2(_16800_),
    .ZN(_05876_));
 AND2_X1 _31006_ (.A1(_05876_),
    .A2(_05870_),
    .ZN(_05877_));
 AND2_X2 _31007_ (.A1(_05746_),
    .A2(_05778_),
    .ZN(_05878_));
 AND2_X1 _31008_ (.A1(_05870_),
    .A2(_05878_),
    .ZN(_05879_));
 AND3_X1 _31009_ (.A1(_05844_),
    .A2(_05749_),
    .A3(_05825_),
    .ZN(_05880_));
 OR4_X1 _31010_ (.A1(_05875_),
    .A2(_05877_),
    .A3(_05879_),
    .A4(_05880_),
    .ZN(_05881_));
 AND2_X1 _31011_ (.A1(_05801_),
    .A2(_05749_),
    .ZN(_05882_));
 CLKBUF_X2 _31012_ (.A(_05882_),
    .Z(_05883_));
 AND2_X1 _31013_ (.A1(_05883_),
    .A2(_05804_),
    .ZN(_05884_));
 BUF_X2 _31014_ (.A(_05883_),
    .Z(_05886_));
 CLKBUF_X2 _31015_ (.A(_05743_),
    .Z(_05887_));
 OAI211_X1 _31016_ (.A(_05886_),
    .B(_05779_),
    .C1(_05763_),
    .C2(_05887_),
    .ZN(_05888_));
 INV_X1 _31017_ (.A(_05866_),
    .ZN(_05889_));
 INV_X1 _31018_ (.A(_05883_),
    .ZN(_05890_));
 OAI21_X1 _31019_ (.A(_05888_),
    .B1(_05889_),
    .B2(_05890_),
    .ZN(_05891_));
 CLKBUF_X2 _31020_ (.A(_05739_),
    .Z(_05892_));
 AND3_X1 _31021_ (.A1(_05886_),
    .A2(_05850_),
    .A3(_05892_),
    .ZN(_05893_));
 NOR4_X1 _31022_ (.A1(_05881_),
    .A2(_05884_),
    .A3(_05891_),
    .A4(_05893_),
    .ZN(_05894_));
 NAND4_X2 _31023_ (.A1(_05798_),
    .A2(_05840_),
    .A3(_05869_),
    .A4(_05894_),
    .ZN(_05895_));
 AND2_X1 _31024_ (.A1(_16805_),
    .A2(_16806_),
    .ZN(_05897_));
 AND2_X1 _31025_ (.A1(_05825_),
    .A2(_05897_),
    .ZN(_05898_));
 CLKBUF_X2 _31026_ (.A(_05898_),
    .Z(_05899_));
 CLKBUF_X2 _31027_ (.A(_05899_),
    .Z(_05900_));
 AND2_X1 _31028_ (.A1(_05773_),
    .A2(_05900_),
    .ZN(_05901_));
 AND2_X1 _31029_ (.A1(_05854_),
    .A2(_05899_),
    .ZN(_05902_));
 AND2_X1 _31030_ (.A1(_05876_),
    .A2(_05899_),
    .ZN(_05903_));
 AND2_X1 _31031_ (.A1(_05899_),
    .A2(_05829_),
    .ZN(_05904_));
 OR4_X1 _31032_ (.A1(_05901_),
    .A2(_05902_),
    .A3(_05903_),
    .A4(_05904_),
    .ZN(_05905_));
 CLKBUF_X2 _31033_ (.A(_05897_),
    .Z(_05906_));
 AND2_X1 _31034_ (.A1(_05906_),
    .A2(_05802_),
    .ZN(_05908_));
 CLKBUF_X2 _31035_ (.A(_05908_),
    .Z(_05909_));
 AND2_X1 _31036_ (.A1(_05834_),
    .A2(_05909_),
    .ZN(_05910_));
 INV_X1 _31037_ (.A(_05910_),
    .ZN(_05911_));
 BUF_X2 _31038_ (.A(_05909_),
    .Z(_05912_));
 AND2_X1 _31039_ (.A1(_05778_),
    .A2(_05745_),
    .ZN(_05913_));
 NAND2_X1 _31040_ (.A1(_05912_),
    .A2(_05913_),
    .ZN(_05914_));
 NAND2_X1 _31041_ (.A1(_05911_),
    .A2(_05914_),
    .ZN(_05915_));
 AND3_X1 _31042_ (.A1(_05899_),
    .A2(_05833_),
    .A3(_05747_),
    .ZN(_05916_));
 AND2_X1 _31043_ (.A1(_05777_),
    .A2(_05762_),
    .ZN(_05917_));
 AND2_X1 _31044_ (.A1(_05899_),
    .A2(_05917_),
    .ZN(_05919_));
 AND3_X1 _31045_ (.A1(_05783_),
    .A2(_05906_),
    .A3(_05825_),
    .ZN(_05920_));
 OR3_X1 _31046_ (.A1(_05916_),
    .A2(_05919_),
    .A3(_05920_),
    .ZN(_05921_));
 INV_X1 _31047_ (.A(_05909_),
    .ZN(_05922_));
 AOI21_X1 _31048_ (.A(_05922_),
    .B1(_05812_),
    .B2(_05873_),
    .ZN(_05923_));
 NOR4_X1 _31049_ (.A1(_05905_),
    .A2(_05915_),
    .A3(_05921_),
    .A4(_05923_),
    .ZN(_05924_));
 AND2_X1 _31050_ (.A1(_05756_),
    .A2(_05906_),
    .ZN(_05925_));
 AND2_X1 _31051_ (.A1(_05925_),
    .A2(_05857_),
    .ZN(_05926_));
 AND2_X1 _31052_ (.A1(_05925_),
    .A2(_05773_),
    .ZN(_05927_));
 NOR2_X1 _31053_ (.A1(_05926_),
    .A2(_05927_),
    .ZN(_05928_));
 AND2_X1 _31054_ (.A1(_05787_),
    .A2(_05767_),
    .ZN(_05930_));
 CLKBUF_X2 _31055_ (.A(_05930_),
    .Z(_05931_));
 AND2_X1 _31056_ (.A1(_05925_),
    .A2(_05931_),
    .ZN(_05932_));
 INV_X1 _31057_ (.A(_05932_),
    .ZN(_05933_));
 OAI211_X1 _31058_ (.A(_05925_),
    .B(_05779_),
    .C1(_05850_),
    .C2(_05781_),
    .ZN(_05934_));
 AND2_X1 _31059_ (.A1(_05933_),
    .A2(_05934_),
    .ZN(_05935_));
 AND3_X1 _31060_ (.A1(_05739_),
    .A2(_05906_),
    .A3(_05748_),
    .ZN(_05936_));
 AND2_X1 _31061_ (.A1(_05762_),
    .A2(_05759_),
    .ZN(_05937_));
 AND2_X1 _31062_ (.A1(_05906_),
    .A2(_05748_),
    .ZN(_05938_));
 BUF_X2 _31063_ (.A(_05938_),
    .Z(_05939_));
 AOI22_X1 _31064_ (.A1(_05936_),
    .A2(_05821_),
    .B1(_05937_),
    .B2(_05939_),
    .ZN(_05941_));
 AND2_X1 _31065_ (.A1(_05789_),
    .A2(_05938_),
    .ZN(_05942_));
 AND2_X1 _31066_ (.A1(_05878_),
    .A2(_05939_),
    .ZN(_05943_));
 AND2_X1 _31067_ (.A1(_05837_),
    .A2(_05938_),
    .ZN(_05944_));
 NOR3_X1 _31068_ (.A1(_05942_),
    .A2(_05943_),
    .A3(_05944_),
    .ZN(_05945_));
 AND4_X1 _31069_ (.A1(_05928_),
    .A2(_05935_),
    .A3(_05941_),
    .A4(_05945_),
    .ZN(_05946_));
 AND2_X1 _31070_ (.A1(_05799_),
    .A2(_16806_),
    .ZN(_05947_));
 CLKBUF_X2 _31071_ (.A(_05947_),
    .Z(_05948_));
 OAI211_X1 _31072_ (.A(_05848_),
    .B(_05948_),
    .C1(_05876_),
    .C2(_05804_),
    .ZN(_05949_));
 AND2_X1 _31073_ (.A1(_05756_),
    .A2(_05947_),
    .ZN(_05950_));
 CLKBUF_X2 _31074_ (.A(_05950_),
    .Z(_05952_));
 INV_X1 _31075_ (.A(_05783_),
    .ZN(_05953_));
 INV_X1 _31076_ (.A(_05917_),
    .ZN(_05954_));
 NAND2_X1 _31077_ (.A1(_05953_),
    .A2(_05954_),
    .ZN(_05955_));
 OAI21_X1 _31078_ (.A(_05952_),
    .B1(_05955_),
    .B2(_05846_),
    .ZN(_05956_));
 AND2_X1 _31079_ (.A1(_05947_),
    .A2(_05748_),
    .ZN(_05957_));
 CLKBUF_X2 _31080_ (.A(_05957_),
    .Z(_05958_));
 AND2_X1 _31081_ (.A1(_05767_),
    .A2(_05758_),
    .ZN(_05959_));
 INV_X1 _31082_ (.A(_05959_),
    .ZN(_05960_));
 INV_X1 _31083_ (.A(_05937_),
    .ZN(_05961_));
 NAND2_X1 _31084_ (.A1(_05960_),
    .A2(_05961_),
    .ZN(_05963_));
 OAI21_X1 _31085_ (.A(_05958_),
    .B1(_05963_),
    .B2(_05855_),
    .ZN(_05964_));
 NAND2_X1 _31086_ (.A1(_05958_),
    .A2(_05789_),
    .ZN(_05965_));
 AND4_X1 _31087_ (.A1(_05949_),
    .A2(_05956_),
    .A3(_05964_),
    .A4(_05965_),
    .ZN(_05966_));
 AND2_X1 _31088_ (.A1(_05947_),
    .A2(_05802_),
    .ZN(_05967_));
 AND2_X1 _31089_ (.A1(_05967_),
    .A2(_05866_),
    .ZN(_05968_));
 AND2_X1 _31090_ (.A1(_05743_),
    .A2(_05777_),
    .ZN(_05969_));
 AND2_X1 _31091_ (.A1(_05967_),
    .A2(_05969_),
    .ZN(_05970_));
 NOR2_X1 _31092_ (.A1(_05968_),
    .A2(_05970_),
    .ZN(_05971_));
 AND2_X1 _31093_ (.A1(_05947_),
    .A2(_05825_),
    .ZN(_05972_));
 CLKBUF_X2 _31094_ (.A(_05972_),
    .Z(_05974_));
 AND2_X1 _31095_ (.A1(_05974_),
    .A2(_05937_),
    .ZN(_05975_));
 INV_X1 _31096_ (.A(_05975_),
    .ZN(_05976_));
 CLKBUF_X2 _31097_ (.A(_05833_),
    .Z(_05977_));
 OAI221_X1 _31098_ (.A(_05974_),
    .B1(_05780_),
    .B2(_05781_),
    .C1(_05779_),
    .C2(_05977_),
    .ZN(_05978_));
 CLKBUF_X2 _31099_ (.A(_05967_),
    .Z(_05979_));
 OAI21_X1 _31100_ (.A(_05979_),
    .B1(_05744_),
    .B2(_05829_),
    .ZN(_05980_));
 AND4_X1 _31101_ (.A1(_05971_),
    .A2(_05976_),
    .A3(_05978_),
    .A4(_05980_),
    .ZN(_05981_));
 NAND4_X2 _31102_ (.A1(_05924_),
    .A2(_05946_),
    .A3(_05966_),
    .A4(_05981_),
    .ZN(_05982_));
 NOR2_X4 _31103_ (.A1(_05895_),
    .A2(_05982_),
    .ZN(_05983_));
 INV_X1 _31104_ (.A(_05983_),
    .ZN(_05985_));
 NOR2_X2 _31105_ (.A1(_16760_),
    .A2(_16759_),
    .ZN(_05986_));
 INV_X2 _31106_ (.A(_05986_),
    .ZN(_05987_));
 AND2_X1 _31107_ (.A1(_16761_),
    .A2(_16762_),
    .ZN(_05988_));
 NAND2_X1 _31108_ (.A1(_05987_),
    .A2(_05988_),
    .ZN(_05989_));
 INV_X1 _31109_ (.A(_05989_),
    .ZN(_05990_));
 AND2_X1 _31110_ (.A1(_16760_),
    .A2(_16759_),
    .ZN(_05991_));
 INV_X1 _31111_ (.A(_05991_),
    .ZN(_05992_));
 NOR2_X2 _31112_ (.A1(_16766_),
    .A2(_16765_),
    .ZN(_05993_));
 NOR2_X2 _31113_ (.A1(_16764_),
    .A2(_16763_),
    .ZN(_05994_));
 AND2_X2 _31114_ (.A1(_05993_),
    .A2(_05994_),
    .ZN(_05996_));
 BUF_X2 _31115_ (.A(_05996_),
    .Z(_05997_));
 NAND3_X1 _31116_ (.A1(_05990_),
    .A2(_05992_),
    .A3(_05997_),
    .ZN(_05998_));
 NOR2_X2 _31117_ (.A1(_16761_),
    .A2(_16762_),
    .ZN(_05999_));
 AND2_X2 _31118_ (.A1(_05999_),
    .A2(_16760_),
    .ZN(_06000_));
 NAND2_X1 _31119_ (.A1(_05996_),
    .A2(_06000_),
    .ZN(_06001_));
 INV_X1 _31120_ (.A(_16761_),
    .ZN(_06002_));
 NOR2_X1 _31121_ (.A1(_06002_),
    .A2(_16762_),
    .ZN(_06003_));
 CLKBUF_X2 _31122_ (.A(_06003_),
    .Z(_06004_));
 CLKBUF_X2 _31123_ (.A(_06004_),
    .Z(_06005_));
 CLKBUF_X2 _31124_ (.A(_06005_),
    .Z(_06007_));
 BUF_X2 _31125_ (.A(_16760_),
    .Z(_06008_));
 CLKBUF_X2 _31126_ (.A(_16759_),
    .Z(_06009_));
 OAI211_X1 _31127_ (.A(_05997_),
    .B(_06007_),
    .C1(_06008_),
    .C2(_06009_),
    .ZN(_06010_));
 INV_X1 _31128_ (.A(_16762_),
    .ZN(_06011_));
 NOR2_X2 _31129_ (.A1(_06011_),
    .A2(_16761_),
    .ZN(_06012_));
 CLKBUF_X2 _31130_ (.A(_06012_),
    .Z(_06013_));
 CLKBUF_X2 _31131_ (.A(_06013_),
    .Z(_06014_));
 OAI211_X1 _31132_ (.A(_05997_),
    .B(_06014_),
    .C1(_06008_),
    .C2(_06009_),
    .ZN(_06015_));
 AND4_X1 _31133_ (.A1(_05998_),
    .A2(_06001_),
    .A3(_06010_),
    .A4(_06015_),
    .ZN(_06016_));
 NAND2_X1 _31134_ (.A1(_05992_),
    .A2(_06004_),
    .ZN(_06018_));
 INV_X1 _31135_ (.A(_06018_),
    .ZN(_06019_));
 INV_X1 _31136_ (.A(_16764_),
    .ZN(_06020_));
 AND2_X1 _31137_ (.A1(_06020_),
    .A2(_16763_),
    .ZN(_06021_));
 AND2_X1 _31138_ (.A1(_06021_),
    .A2(_05993_),
    .ZN(_06022_));
 CLKBUF_X2 _31139_ (.A(_06022_),
    .Z(_06023_));
 AND3_X1 _31140_ (.A1(_06019_),
    .A2(_05987_),
    .A3(_06023_),
    .ZN(_06024_));
 INV_X1 _31141_ (.A(_06012_),
    .ZN(_06025_));
 INV_X1 _31142_ (.A(_16759_),
    .ZN(_06026_));
 NOR2_X2 _31143_ (.A1(_06026_),
    .A2(_16760_),
    .ZN(_06027_));
 OR2_X1 _31144_ (.A1(_06025_),
    .A2(_06027_),
    .ZN(_06029_));
 INV_X1 _31145_ (.A(_16760_),
    .ZN(_06030_));
 NOR2_X1 _31146_ (.A1(_06030_),
    .A2(_16759_),
    .ZN(_06031_));
 CLKBUF_X2 _31147_ (.A(_06031_),
    .Z(_06032_));
 NOR2_X1 _31148_ (.A1(_06029_),
    .A2(_06032_),
    .ZN(_06033_));
 AND2_X1 _31149_ (.A1(_06033_),
    .A2(_06023_),
    .ZN(_06034_));
 BUF_X2 _31150_ (.A(_06023_),
    .Z(_06035_));
 AOI211_X1 _31151_ (.A(_06024_),
    .B(_06034_),
    .C1(_06000_),
    .C2(_06035_),
    .ZN(_06036_));
 NOR2_X2 _31152_ (.A1(_06020_),
    .A2(_16763_),
    .ZN(_06037_));
 AND2_X2 _31153_ (.A1(_06037_),
    .A2(_05993_),
    .ZN(_06038_));
 INV_X1 _31154_ (.A(_06038_),
    .ZN(_06040_));
 NOR2_X1 _31155_ (.A1(_06018_),
    .A2(_05986_),
    .ZN(_06041_));
 INV_X1 _31156_ (.A(_06041_),
    .ZN(_06042_));
 CLKBUF_X2 _31157_ (.A(_05999_),
    .Z(_06043_));
 BUF_X2 _31158_ (.A(_06030_),
    .Z(_06044_));
 CLKBUF_X2 _31159_ (.A(_06026_),
    .Z(_06045_));
 OAI21_X1 _31160_ (.A(_06043_),
    .B1(_06044_),
    .B2(_06045_),
    .ZN(_06046_));
 AOI21_X1 _31161_ (.A(_06040_),
    .B1(_06042_),
    .B2(_06046_),
    .ZN(_06047_));
 AND2_X1 _31162_ (.A1(_05988_),
    .A2(_16760_),
    .ZN(_06048_));
 BUF_X2 _31163_ (.A(_06048_),
    .Z(_06049_));
 AND2_X1 _31164_ (.A1(_06038_),
    .A2(_06049_),
    .ZN(_06051_));
 AND2_X2 _31165_ (.A1(_05988_),
    .A2(_05986_),
    .ZN(_06052_));
 AND3_X1 _31166_ (.A1(_06052_),
    .A2(_05993_),
    .A3(_06037_),
    .ZN(_06053_));
 NAND2_X1 _31167_ (.A1(_05987_),
    .A2(_06013_),
    .ZN(_06054_));
 INV_X1 _31168_ (.A(_06054_),
    .ZN(_06055_));
 AND2_X1 _31169_ (.A1(_06055_),
    .A2(_06038_),
    .ZN(_06056_));
 NOR4_X1 _31170_ (.A1(_06047_),
    .A2(_06051_),
    .A3(_06053_),
    .A4(_06056_),
    .ZN(_06057_));
 CLKBUF_X2 _31171_ (.A(_05988_),
    .Z(_06058_));
 BUF_X2 _31172_ (.A(_06058_),
    .Z(_06059_));
 INV_X1 _31173_ (.A(_06059_),
    .ZN(_06060_));
 AND2_X1 _31174_ (.A1(_16764_),
    .A2(_16763_),
    .ZN(_06062_));
 AND2_X2 _31175_ (.A1(_06062_),
    .A2(_05993_),
    .ZN(_06063_));
 INV_X1 _31176_ (.A(_06063_),
    .ZN(_06064_));
 CLKBUF_X2 _31177_ (.A(_06045_),
    .Z(_06065_));
 AOI211_X1 _31178_ (.A(_06060_),
    .B(_06064_),
    .C1(_06008_),
    .C2(_06065_),
    .ZN(_06066_));
 NAND2_X1 _31179_ (.A1(_05987_),
    .A2(_05999_),
    .ZN(_06067_));
 NOR2_X1 _31180_ (.A1(_06064_),
    .A2(_06067_),
    .ZN(_06068_));
 AND2_X1 _31181_ (.A1(_06012_),
    .A2(_05986_),
    .ZN(_06069_));
 AND2_X1 _31182_ (.A1(_06069_),
    .A2(_06063_),
    .ZN(_06070_));
 AND3_X1 _31183_ (.A1(_06063_),
    .A2(_06005_),
    .A3(_06032_),
    .ZN(_06071_));
 NOR4_X1 _31184_ (.A1(_06066_),
    .A2(_06068_),
    .A3(_06070_),
    .A4(_06071_),
    .ZN(_06073_));
 AND4_X1 _31185_ (.A1(_06016_),
    .A2(_06036_),
    .A3(_06057_),
    .A4(_06073_),
    .ZN(_06074_));
 AND2_X1 _31186_ (.A1(_06027_),
    .A2(_06043_),
    .ZN(_06075_));
 CLKBUF_X2 _31187_ (.A(_06075_),
    .Z(_06076_));
 AND2_X1 _31188_ (.A1(_16766_),
    .A2(_16765_),
    .ZN(_06077_));
 AND2_X2 _31189_ (.A1(_06077_),
    .A2(_06062_),
    .ZN(_06078_));
 AND2_X1 _31190_ (.A1(_06076_),
    .A2(_06078_),
    .ZN(_06079_));
 AND2_X1 _31191_ (.A1(_06004_),
    .A2(_05986_),
    .ZN(_06080_));
 AND2_X1 _31192_ (.A1(_06080_),
    .A2(_06078_),
    .ZN(_06081_));
 CLKBUF_X2 _31193_ (.A(_06078_),
    .Z(_06082_));
 AOI211_X1 _31194_ (.A(_06079_),
    .B(_06081_),
    .C1(_06000_),
    .C2(_06082_),
    .ZN(_06084_));
 AND2_X1 _31195_ (.A1(_06031_),
    .A2(_05988_),
    .ZN(_06085_));
 CLKBUF_X2 _31196_ (.A(_06085_),
    .Z(_06086_));
 NAND2_X1 _31197_ (.A1(_06086_),
    .A2(_06082_),
    .ZN(_06087_));
 INV_X1 _31198_ (.A(_06078_),
    .ZN(_06088_));
 OAI211_X1 _31199_ (.A(_06084_),
    .B(_06087_),
    .C1(_06025_),
    .C2(_06088_),
    .ZN(_06089_));
 AND2_X1 _31200_ (.A1(_06021_),
    .A2(_06077_),
    .ZN(_06090_));
 AND2_X2 _31201_ (.A1(_06031_),
    .A2(_06012_),
    .ZN(_06091_));
 AND2_X1 _31202_ (.A1(_06090_),
    .A2(_06091_),
    .ZN(_06092_));
 AND2_X1 _31203_ (.A1(_06012_),
    .A2(_05991_),
    .ZN(_06093_));
 CLKBUF_X2 _31204_ (.A(_06093_),
    .Z(_06095_));
 AND2_X1 _31205_ (.A1(_06090_),
    .A2(_06095_),
    .ZN(_06096_));
 BUF_X2 _31206_ (.A(_06090_),
    .Z(_06097_));
 NAND2_X2 _31207_ (.A1(_06012_),
    .A2(_06030_),
    .ZN(_06098_));
 INV_X2 _31208_ (.A(_06098_),
    .ZN(_06099_));
 AOI211_X1 _31209_ (.A(_06092_),
    .B(_06096_),
    .C1(_06097_),
    .C2(_06099_),
    .ZN(_06100_));
 AND2_X2 _31210_ (.A1(_06004_),
    .A2(_06027_),
    .ZN(_06101_));
 AND2_X1 _31211_ (.A1(_06031_),
    .A2(_05999_),
    .ZN(_06102_));
 CLKBUF_X2 _31212_ (.A(_06102_),
    .Z(_06103_));
 OAI21_X1 _31213_ (.A(_06097_),
    .B1(_06101_),
    .B2(_06103_),
    .ZN(_06104_));
 AND2_X1 _31214_ (.A1(_06027_),
    .A2(_05988_),
    .ZN(_06106_));
 BUF_X2 _31215_ (.A(_06106_),
    .Z(_06107_));
 OAI21_X1 _31216_ (.A(_06097_),
    .B1(_06107_),
    .B2(_06086_),
    .ZN(_06108_));
 NAND3_X1 _31217_ (.A1(_06100_),
    .A2(_06104_),
    .A3(_06108_),
    .ZN(_06109_));
 AND2_X2 _31218_ (.A1(_06077_),
    .A2(_05994_),
    .ZN(_06110_));
 BUF_X2 _31219_ (.A(_06110_),
    .Z(_06111_));
 OAI211_X1 _31220_ (.A(_06111_),
    .B(_06059_),
    .C1(_06044_),
    .C2(_06065_),
    .ZN(_06112_));
 NAND2_X1 _31221_ (.A1(_06103_),
    .A2(_06111_),
    .ZN(_06113_));
 AND2_X1 _31222_ (.A1(_06013_),
    .A2(_06009_),
    .ZN(_06114_));
 INV_X1 _31223_ (.A(_06114_),
    .ZN(_06115_));
 INV_X1 _31224_ (.A(_06110_),
    .ZN(_06117_));
 OAI211_X1 _31225_ (.A(_06112_),
    .B(_06113_),
    .C1(_06115_),
    .C2(_06117_),
    .ZN(_06118_));
 AND2_X1 _31226_ (.A1(_06037_),
    .A2(_06077_),
    .ZN(_06119_));
 INV_X1 _31227_ (.A(_06119_),
    .ZN(_06120_));
 NOR2_X1 _31228_ (.A1(_06029_),
    .A2(_06120_),
    .ZN(_06121_));
 CLKBUF_X2 _31229_ (.A(_06119_),
    .Z(_06122_));
 INV_X1 _31230_ (.A(_06043_),
    .ZN(_06123_));
 NOR2_X1 _31231_ (.A1(_06123_),
    .A2(_06027_),
    .ZN(_06124_));
 INV_X1 _31232_ (.A(_06031_),
    .ZN(_06125_));
 AND3_X1 _31233_ (.A1(_06122_),
    .A2(_06124_),
    .A3(_06125_),
    .ZN(_06126_));
 AND2_X1 _31234_ (.A1(_06004_),
    .A2(_06030_),
    .ZN(_06128_));
 AND2_X1 _31235_ (.A1(_06128_),
    .A2(_06119_),
    .ZN(_06129_));
 AND2_X1 _31236_ (.A1(_06058_),
    .A2(_16759_),
    .ZN(_06130_));
 AND2_X1 _31237_ (.A1(_06119_),
    .A2(_06130_),
    .ZN(_06131_));
 OR4_X1 _31238_ (.A1(_06121_),
    .A2(_06126_),
    .A3(_06129_),
    .A4(_06131_),
    .ZN(_06132_));
 NOR4_X1 _31239_ (.A1(_06089_),
    .A2(_06109_),
    .A3(_06118_),
    .A4(_06132_),
    .ZN(_06133_));
 INV_X1 _31240_ (.A(_16766_),
    .ZN(_06134_));
 AND2_X1 _31241_ (.A1(_06134_),
    .A2(_16765_),
    .ZN(_06135_));
 AND2_X1 _31242_ (.A1(_06135_),
    .A2(_05994_),
    .ZN(_06136_));
 BUF_X2 _31243_ (.A(_06136_),
    .Z(_06137_));
 AND2_X1 _31244_ (.A1(_06137_),
    .A2(_06080_),
    .ZN(_06139_));
 INV_X1 _31245_ (.A(_06137_),
    .ZN(_06140_));
 AOI22_X1 _31246_ (.A1(_05992_),
    .A2(_06059_),
    .B1(_06013_),
    .B2(_06009_),
    .ZN(_06141_));
 NOR2_X1 _31247_ (.A1(_06140_),
    .A2(_06141_),
    .ZN(_06142_));
 AND2_X2 _31248_ (.A1(_05999_),
    .A2(_06030_),
    .ZN(_06143_));
 AOI211_X1 _31249_ (.A(_06139_),
    .B(_06142_),
    .C1(_06143_),
    .C2(_06137_),
    .ZN(_06144_));
 AND2_X2 _31250_ (.A1(_06135_),
    .A2(_06037_),
    .ZN(_06145_));
 AND2_X2 _31251_ (.A1(_06004_),
    .A2(_06031_),
    .ZN(_06146_));
 AND2_X1 _31252_ (.A1(_06145_),
    .A2(_06146_),
    .ZN(_06147_));
 INV_X1 _31253_ (.A(_06147_),
    .ZN(_06148_));
 BUF_X2 _31254_ (.A(_05991_),
    .Z(_06150_));
 AND2_X2 _31255_ (.A1(_06004_),
    .A2(_06150_),
    .ZN(_06151_));
 NAND2_X1 _31256_ (.A1(_06145_),
    .A2(_06151_),
    .ZN(_06152_));
 CLKBUF_X2 _31257_ (.A(_06145_),
    .Z(_06153_));
 NAND2_X1 _31258_ (.A1(_06153_),
    .A2(_06128_),
    .ZN(_06154_));
 NAND3_X1 _31259_ (.A1(_06148_),
    .A2(_06152_),
    .A3(_06154_),
    .ZN(_06155_));
 AND2_X1 _31260_ (.A1(_06145_),
    .A2(_06076_),
    .ZN(_06156_));
 NAND2_X1 _31261_ (.A1(_06145_),
    .A2(_06085_),
    .ZN(_06157_));
 CLKBUF_X2 _31262_ (.A(_06135_),
    .Z(_06158_));
 NAND4_X1 _31263_ (.A1(_06158_),
    .A2(_06013_),
    .A3(_06037_),
    .A4(_06150_),
    .ZN(_06159_));
 INV_X1 _31264_ (.A(_06145_),
    .ZN(_06161_));
 OAI211_X1 _31265_ (.A(_06157_),
    .B(_06159_),
    .C1(_06161_),
    .C2(_06098_),
    .ZN(_06162_));
 AND2_X1 _31266_ (.A1(_05991_),
    .A2(_05999_),
    .ZN(_06163_));
 AND2_X1 _31267_ (.A1(_06145_),
    .A2(_06163_),
    .ZN(_06164_));
 NOR4_X1 _31268_ (.A1(_06155_),
    .A2(_06156_),
    .A3(_06162_),
    .A4(_06164_),
    .ZN(_06165_));
 AND2_X1 _31269_ (.A1(_06135_),
    .A2(_06021_),
    .ZN(_06166_));
 BUF_X2 _31270_ (.A(_06166_),
    .Z(_06167_));
 AND2_X2 _31271_ (.A1(_06004_),
    .A2(_16760_),
    .ZN(_06168_));
 AND2_X1 _31272_ (.A1(_06167_),
    .A2(_06168_),
    .ZN(_06169_));
 AND2_X2 _31273_ (.A1(_06150_),
    .A2(_05988_),
    .ZN(_06170_));
 CLKBUF_X2 _31274_ (.A(_06021_),
    .Z(_06172_));
 NAND3_X1 _31275_ (.A1(_06170_),
    .A2(_06172_),
    .A3(_06158_),
    .ZN(_06173_));
 INV_X1 _31276_ (.A(_06166_),
    .ZN(_06174_));
 OAI21_X1 _31277_ (.A(_06173_),
    .B1(_06174_),
    .B2(_06115_),
    .ZN(_06175_));
 OAI21_X1 _31278_ (.A(_06043_),
    .B1(_06044_),
    .B2(_16759_),
    .ZN(_06176_));
 INV_X1 _31279_ (.A(_06176_),
    .ZN(_06177_));
 AOI211_X1 _31280_ (.A(_06169_),
    .B(_06175_),
    .C1(_06167_),
    .C2(_06177_),
    .ZN(_06178_));
 AND2_X1 _31281_ (.A1(_06135_),
    .A2(_06062_),
    .ZN(_06179_));
 BUF_X2 _31282_ (.A(_06179_),
    .Z(_06180_));
 OAI21_X1 _31283_ (.A(_06180_),
    .B1(_06107_),
    .B2(_06085_),
    .ZN(_06181_));
 CLKBUF_X2 _31284_ (.A(_06062_),
    .Z(_06183_));
 NAND3_X1 _31285_ (.A1(_06095_),
    .A2(_06158_),
    .A3(_06183_),
    .ZN(_06184_));
 NAND2_X1 _31286_ (.A1(_06181_),
    .A2(_06184_),
    .ZN(_06185_));
 INV_X1 _31287_ (.A(_06185_),
    .ZN(_06186_));
 NAND2_X1 _31288_ (.A1(_06180_),
    .A2(_06163_),
    .ZN(_06187_));
 AND2_X1 _31289_ (.A1(_06003_),
    .A2(_16759_),
    .ZN(_06188_));
 NAND2_X1 _31290_ (.A1(_06180_),
    .A2(_06188_),
    .ZN(_06189_));
 AND2_X1 _31291_ (.A1(_05999_),
    .A2(_05986_),
    .ZN(_06190_));
 OAI21_X1 _31292_ (.A(_06180_),
    .B1(_06076_),
    .B2(_06190_),
    .ZN(_06191_));
 AND4_X1 _31293_ (.A1(_06186_),
    .A2(_06187_),
    .A3(_06189_),
    .A4(_06191_),
    .ZN(_06192_));
 AND4_X1 _31294_ (.A1(_06144_),
    .A2(_06165_),
    .A3(_06178_),
    .A4(_06192_),
    .ZN(_06194_));
 NOR2_X1 _31295_ (.A1(_06134_),
    .A2(_16765_),
    .ZN(_06195_));
 AND2_X1 _31296_ (.A1(_06021_),
    .A2(_06195_),
    .ZN(_06196_));
 BUF_X2 _31297_ (.A(_06196_),
    .Z(_06197_));
 BUF_X2 _31298_ (.A(_06027_),
    .Z(_06198_));
 OAI21_X1 _31299_ (.A(_06043_),
    .B1(_06198_),
    .B2(_06032_),
    .ZN(_06199_));
 INV_X1 _31300_ (.A(_06199_),
    .ZN(_06200_));
 OAI21_X1 _31301_ (.A(_06197_),
    .B1(_06200_),
    .B2(_06049_),
    .ZN(_06201_));
 AND2_X2 _31302_ (.A1(_06195_),
    .A2(_06183_),
    .ZN(_06202_));
 OAI21_X1 _31303_ (.A(_06202_),
    .B1(_06190_),
    .B2(_06000_),
    .ZN(_06203_));
 NAND2_X1 _31304_ (.A1(_06125_),
    .A2(_06005_),
    .ZN(_06205_));
 INV_X1 _31305_ (.A(_06202_),
    .ZN(_06206_));
 OAI21_X1 _31306_ (.A(_06203_),
    .B1(_06205_),
    .B2(_06206_),
    .ZN(_06207_));
 AND2_X1 _31307_ (.A1(_06037_),
    .A2(_06195_),
    .ZN(_06208_));
 CLKBUF_X2 _31308_ (.A(_06208_),
    .Z(_06209_));
 CLKBUF_X2 _31309_ (.A(_06209_),
    .Z(_06210_));
 AND2_X1 _31310_ (.A1(_06058_),
    .A2(_06030_),
    .ZN(_06211_));
 OAI21_X1 _31311_ (.A(_06210_),
    .B1(_06170_),
    .B2(_06211_),
    .ZN(_06212_));
 CLKBUF_X2 _31312_ (.A(_06195_),
    .Z(_06213_));
 NAND4_X1 _31313_ (.A1(_06198_),
    .A2(_06014_),
    .A3(_06037_),
    .A4(_06213_),
    .ZN(_06214_));
 NAND2_X1 _31314_ (.A1(_06212_),
    .A2(_06214_),
    .ZN(_06216_));
 AND2_X1 _31315_ (.A1(_06209_),
    .A2(_06080_),
    .ZN(_06217_));
 AND3_X1 _31316_ (.A1(_06052_),
    .A2(_06213_),
    .A3(_06183_),
    .ZN(_06218_));
 NOR4_X1 _31317_ (.A1(_06207_),
    .A2(_06216_),
    .A3(_06217_),
    .A4(_06218_),
    .ZN(_06219_));
 AND4_X1 _31318_ (.A1(_06005_),
    .A2(_06213_),
    .A3(_06150_),
    .A4(_05994_),
    .ZN(_06220_));
 AND2_X2 _31319_ (.A1(_06195_),
    .A2(_05994_),
    .ZN(_06221_));
 AND2_X1 _31320_ (.A1(_06128_),
    .A2(_06221_),
    .ZN(_06222_));
 AND2_X1 _31321_ (.A1(_06043_),
    .A2(_06045_),
    .ZN(_06223_));
 BUF_X2 _31322_ (.A(_06221_),
    .Z(_06224_));
 AOI211_X1 _31323_ (.A(_06220_),
    .B(_06222_),
    .C1(_06223_),
    .C2(_06224_),
    .ZN(_06225_));
 OAI21_X1 _31324_ (.A(_06224_),
    .B1(_05990_),
    .B2(_06114_),
    .ZN(_06227_));
 AND4_X1 _31325_ (.A1(_06201_),
    .A2(_06219_),
    .A3(_06225_),
    .A4(_06227_),
    .ZN(_06228_));
 NAND4_X1 _31326_ (.A1(_06074_),
    .A2(_06133_),
    .A3(_06194_),
    .A4(_06228_),
    .ZN(_06229_));
 OAI21_X1 _31327_ (.A(_06011_),
    .B1(_05987_),
    .B2(_16761_),
    .ZN(_06230_));
 AND3_X1 _31328_ (.A1(_05993_),
    .A2(_05994_),
    .A3(_06011_),
    .ZN(_06231_));
 AND2_X1 _31329_ (.A1(_06230_),
    .A2(_06231_),
    .ZN(_06232_));
 NOR2_X2 _31330_ (.A1(_06229_),
    .A2(_06232_),
    .ZN(_06233_));
 XNOR2_X1 _31331_ (.A(_05985_),
    .B(_06233_),
    .ZN(_06234_));
 XNOR2_X1 _31332_ (.A(_05736_),
    .B(_06234_),
    .ZN(_06235_));
 MUX2_X1 _31333_ (.A(_05121_),
    .B(_06235_),
    .S(_05069_),
    .Z(_00700_));
 MUX2_X1 _31334_ (.A(_17058_),
    .B(_16930_),
    .S(_05119_),
    .Z(_00855_));
 MUX2_X1 _31335_ (.A(_17059_),
    .B(_16931_),
    .S(_05119_),
    .Z(_00856_));
 MUX2_X1 _31336_ (.A(_17060_),
    .B(_16932_),
    .S(_05119_),
    .Z(_00857_));
 MUX2_X1 _31337_ (.A(_17061_),
    .B(_16933_),
    .S(_05119_),
    .Z(_00858_));
 MUX2_X1 _31338_ (.A(_16936_),
    .B(_16808_),
    .S(_05119_),
    .Z(_00733_));
 BUF_X2 _31339_ (.A(_05104_),
    .Z(_06237_));
 MUX2_X1 _31340_ (.A(_16937_),
    .B(_16809_),
    .S(_06237_),
    .Z(_00734_));
 MUX2_X1 _31341_ (.A(_16938_),
    .B(_16810_),
    .S(_06237_),
    .Z(_00735_));
 MUX2_X1 _31342_ (.A(_16939_),
    .B(_16811_),
    .S(_06237_),
    .Z(_00736_));
 MUX2_X1 _31343_ (.A(_16940_),
    .B(_16812_),
    .S(_06237_),
    .Z(_00737_));
 MUX2_X1 _31344_ (.A(_16941_),
    .B(_16813_),
    .S(_06237_),
    .Z(_00738_));
 XOR2_X1 _31345_ (.A(_17110_),
    .B(_17059_),
    .Z(_06239_));
 AND2_X1 _31346_ (.A1(_05524_),
    .A2(_05590_),
    .ZN(_06240_));
 OAI21_X1 _31347_ (.A(_05541_),
    .B1(_06240_),
    .B2(_05616_),
    .ZN(_06241_));
 CLKBUF_X2 _31348_ (.A(_05529_),
    .Z(_06242_));
 NAND3_X1 _31349_ (.A1(_05508_),
    .A2(_06242_),
    .A3(_05486_),
    .ZN(_06243_));
 INV_X1 _31350_ (.A(_05605_),
    .ZN(_06244_));
 INV_X1 _31351_ (.A(_05530_),
    .ZN(_06245_));
 OAI211_X1 _31352_ (.A(_06241_),
    .B(_06243_),
    .C1(_06244_),
    .C2(_06245_),
    .ZN(_06246_));
 INV_X1 _31353_ (.A(_05631_),
    .ZN(_06247_));
 INV_X1 _31354_ (.A(_05704_),
    .ZN(_06249_));
 AOI21_X1 _31355_ (.A(_05563_),
    .B1(_06247_),
    .B2(_06249_),
    .ZN(_06250_));
 BUF_X2 _31356_ (.A(_05562_),
    .Z(_06251_));
 AOI211_X1 _31357_ (.A(_05576_),
    .B(_06250_),
    .C1(_05605_),
    .C2(_06251_),
    .ZN(_06252_));
 NAND2_X1 _31358_ (.A1(_05537_),
    .A2(_05524_),
    .ZN(_06253_));
 INV_X1 _31359_ (.A(_06253_),
    .ZN(_06254_));
 NAND2_X1 _31360_ (.A1(_06254_),
    .A2(_05547_),
    .ZN(_06255_));
 NAND4_X1 _31361_ (.A1(_05666_),
    .A2(_05715_),
    .A3(_05506_),
    .A4(_05596_),
    .ZN(_06256_));
 INV_X1 _31362_ (.A(_05568_),
    .ZN(_06257_));
 OAI21_X1 _31363_ (.A(_06251_),
    .B1(_06257_),
    .B2(_05624_),
    .ZN(_06258_));
 NAND4_X1 _31364_ (.A1(_06252_),
    .A2(_06255_),
    .A3(_06256_),
    .A4(_06258_),
    .ZN(_06260_));
 INV_X1 _31365_ (.A(_05516_),
    .ZN(_06261_));
 AOI21_X1 _31366_ (.A(_05510_),
    .B1(_06261_),
    .B2(_06253_),
    .ZN(_06262_));
 INV_X1 _31367_ (.A(_05492_),
    .ZN(_06263_));
 AOI21_X1 _31368_ (.A(_05510_),
    .B1(_05509_),
    .B2(_06263_),
    .ZN(_06264_));
 NOR4_X1 _31369_ (.A1(_06246_),
    .A2(_06260_),
    .A3(_06262_),
    .A4(_06264_),
    .ZN(_06265_));
 BUF_X2 _31370_ (.A(_05609_),
    .Z(_06266_));
 AND2_X2 _31371_ (.A1(_05524_),
    .A2(_05535_),
    .ZN(_06267_));
 AND2_X2 _31372_ (.A1(_05514_),
    .A2(_05531_),
    .ZN(_06268_));
 OAI21_X1 _31373_ (.A(_06266_),
    .B1(_06267_),
    .B2(_06268_),
    .ZN(_06269_));
 NOR2_X2 _31374_ (.A1(_06263_),
    .A2(_05495_),
    .ZN(_06271_));
 BUF_X2 _31375_ (.A(_06242_),
    .Z(_06272_));
 CLKBUF_X2 _31376_ (.A(_05581_),
    .Z(_06273_));
 NAND4_X1 _31377_ (.A1(_06271_),
    .A2(_06272_),
    .A3(_05666_),
    .A4(_06273_),
    .ZN(_06274_));
 AND2_X1 _31378_ (.A1(_05504_),
    .A2(_05496_),
    .ZN(_06275_));
 NAND2_X1 _31379_ (.A1(_06266_),
    .A2(_06275_),
    .ZN(_06276_));
 NAND2_X1 _31380_ (.A1(_06266_),
    .A2(_05705_),
    .ZN(_06277_));
 NAND4_X1 _31381_ (.A1(_06269_),
    .A2(_06274_),
    .A3(_06276_),
    .A4(_06277_),
    .ZN(_06278_));
 OAI21_X1 _31382_ (.A(_05606_),
    .B1(_05605_),
    .B2(_05703_),
    .ZN(_06279_));
 OAI21_X1 _31383_ (.A(_05606_),
    .B1(_05646_),
    .B2(_05543_),
    .ZN(_06280_));
 INV_X1 _31384_ (.A(_06240_),
    .ZN(_06282_));
 OAI211_X1 _31385_ (.A(_06279_),
    .B(_06280_),
    .C1(_05598_),
    .C2(_06282_),
    .ZN(_06283_));
 OAI21_X1 _31386_ (.A(_05626_),
    .B1(_05674_),
    .B2(_05601_),
    .ZN(_06284_));
 CLKBUF_X2 _31387_ (.A(_05505_),
    .Z(_06285_));
 NAND4_X1 _31388_ (.A1(_05626_),
    .A2(_06285_),
    .A3(_05537_),
    .A4(_05532_),
    .ZN(_06286_));
 INV_X1 _31389_ (.A(_05625_),
    .ZN(_06287_));
 OAI211_X1 _31390_ (.A(_06284_),
    .B(_06286_),
    .C1(_06287_),
    .C2(_05655_),
    .ZN(_06288_));
 OAI211_X1 _31391_ (.A(_05583_),
    .B(_05589_),
    .C1(_05713_),
    .C2(_05499_),
    .ZN(_06289_));
 OAI21_X1 _31392_ (.A(_05582_),
    .B1(_05508_),
    .B2(_05705_),
    .ZN(_06290_));
 BUF_X2 _31393_ (.A(_05524_),
    .Z(_06291_));
 NAND3_X1 _31394_ (.A1(_05583_),
    .A2(_06291_),
    .A3(_05537_),
    .ZN(_06293_));
 NAND4_X1 _31395_ (.A1(_06273_),
    .A2(_05611_),
    .A3(_05715_),
    .A4(_05716_),
    .ZN(_06294_));
 NAND4_X1 _31396_ (.A1(_06289_),
    .A2(_06290_),
    .A3(_06293_),
    .A4(_06294_),
    .ZN(_06295_));
 NOR4_X1 _31397_ (.A1(_06278_),
    .A2(_06283_),
    .A3(_06288_),
    .A4(_06295_),
    .ZN(_06296_));
 AND2_X1 _31398_ (.A1(_05642_),
    .A2(_05644_),
    .ZN(_06297_));
 AND2_X1 _31399_ (.A1(_05642_),
    .A2(_05704_),
    .ZN(_06298_));
 AND2_X1 _31400_ (.A1(_05642_),
    .A2(_05589_),
    .ZN(_06299_));
 AND2_X1 _31401_ (.A1(_05642_),
    .A2(_05690_),
    .ZN(_06300_));
 OR4_X1 _31402_ (.A1(_06297_),
    .A2(_06298_),
    .A3(_06299_),
    .A4(_06300_),
    .ZN(_06301_));
 NAND2_X1 _31403_ (.A1(_05532_),
    .A2(_05504_),
    .ZN(_06302_));
 INV_X1 _31404_ (.A(_06302_),
    .ZN(_06304_));
 AND3_X1 _31405_ (.A1(_06304_),
    .A2(_05651_),
    .A3(_05537_),
    .ZN(_06305_));
 AND2_X1 _31406_ (.A1(_05651_),
    .A2(_05570_),
    .ZN(_06306_));
 AND4_X1 _31407_ (.A1(_05496_),
    .A2(_05637_),
    .A3(_05567_),
    .A4(_05488_),
    .ZN(_06307_));
 OR4_X1 _31408_ (.A1(_05659_),
    .A2(_06305_),
    .A3(_06306_),
    .A4(_06307_),
    .ZN(_06308_));
 CLKBUF_X2 _31409_ (.A(_05561_),
    .Z(_06309_));
 AND4_X1 _31410_ (.A1(_05593_),
    .A2(_05638_),
    .A3(_05567_),
    .A4(_06309_),
    .ZN(_06310_));
 AOI21_X1 _31411_ (.A(_06310_),
    .B1(_05564_),
    .B2(_05670_),
    .ZN(_06311_));
 CLKBUF_X2 _31412_ (.A(_05638_),
    .Z(_06312_));
 NAND4_X1 _31413_ (.A1(_06312_),
    .A2(_05611_),
    .A3(_06285_),
    .A4(_06309_),
    .ZN(_06313_));
 OAI21_X1 _31414_ (.A(_05670_),
    .B1(_05605_),
    .B2(_05701_),
    .ZN(_06315_));
 NAND3_X1 _31415_ (.A1(_06311_),
    .A2(_06313_),
    .A3(_06315_),
    .ZN(_06316_));
 OAI21_X1 _31416_ (.A(_05673_),
    .B1(_05646_),
    .B2(_05543_),
    .ZN(_06317_));
 NAND2_X1 _31417_ (.A1(_05673_),
    .A2(_05699_),
    .ZN(_06318_));
 INV_X1 _31418_ (.A(_05673_),
    .ZN(_06319_));
 OAI211_X1 _31419_ (.A(_06317_),
    .B(_06318_),
    .C1(_05539_),
    .C2(_06319_),
    .ZN(_06320_));
 NOR4_X1 _31420_ (.A1(_06301_),
    .A2(_06308_),
    .A3(_06316_),
    .A4(_06320_),
    .ZN(_06321_));
 NAND3_X1 _31421_ (.A1(_05699_),
    .A2(_06272_),
    .A3(_05714_),
    .ZN(_06322_));
 NAND3_X1 _31422_ (.A1(_05521_),
    .A2(_06272_),
    .A3(_05714_),
    .ZN(_06323_));
 INV_X1 _31423_ (.A(_05696_),
    .ZN(_06324_));
 OAI211_X1 _31424_ (.A(_06322_),
    .B(_06323_),
    .C1(_06324_),
    .C2(_05602_),
    .ZN(_06326_));
 NAND3_X1 _31425_ (.A1(_05570_),
    .A2(_06272_),
    .A3(_05714_),
    .ZN(_06327_));
 NAND4_X1 _31426_ (.A1(_06242_),
    .A2(_06285_),
    .A3(_05496_),
    .A4(_05679_),
    .ZN(_06328_));
 INV_X1 _31427_ (.A(_05557_),
    .ZN(_06329_));
 OAI211_X1 _31428_ (.A(_06327_),
    .B(_06328_),
    .C1(_06324_),
    .C2(_06329_),
    .ZN(_06330_));
 NAND2_X1 _31429_ (.A1(_05633_),
    .A2(_05710_),
    .ZN(_06331_));
 NAND2_X1 _31430_ (.A1(_05710_),
    .A2(_05557_),
    .ZN(_06332_));
 OAI211_X1 _31431_ (.A(_06331_),
    .B(_06332_),
    .C1(_05648_),
    .C2(_05718_),
    .ZN(_06333_));
 OAI21_X1 _31432_ (.A(_05710_),
    .B1(_05619_),
    .B2(_06268_),
    .ZN(_06334_));
 INV_X1 _31433_ (.A(_05624_),
    .ZN(_06335_));
 OAI21_X1 _31434_ (.A(_06334_),
    .B1(_06335_),
    .B2(_05718_),
    .ZN(_06337_));
 NOR4_X1 _31435_ (.A1(_06326_),
    .A2(_06330_),
    .A3(_06333_),
    .A4(_06337_),
    .ZN(_06338_));
 AND3_X1 _31436_ (.A1(_06271_),
    .A2(_05681_),
    .A3(_05664_),
    .ZN(_06339_));
 NAND2_X1 _31437_ (.A1(_05681_),
    .A2(_05705_),
    .ZN(_06340_));
 INV_X1 _31438_ (.A(_06275_),
    .ZN(_06341_));
 OAI21_X1 _31439_ (.A(_06340_),
    .B1(_06341_),
    .B2(_05682_),
    .ZN(_06342_));
 BUF_X2 _31440_ (.A(_05681_),
    .Z(_06343_));
 AOI211_X1 _31441_ (.A(_06339_),
    .B(_06342_),
    .C1(_05564_),
    .C2(_06343_),
    .ZN(_06344_));
 OAI211_X1 _31442_ (.A(_05722_),
    .B(_06291_),
    .C1(_05711_),
    .C2(_05593_),
    .ZN(_06345_));
 BUF_X2 _31443_ (.A(_05558_),
    .Z(_06346_));
 OAI21_X1 _31444_ (.A(_05722_),
    .B1(_05633_),
    .B2(_06346_),
    .ZN(_06348_));
 AND4_X1 _31445_ (.A1(_06338_),
    .A2(_06344_),
    .A3(_06345_),
    .A4(_06348_),
    .ZN(_06349_));
 NAND4_X1 _31446_ (.A1(_06265_),
    .A2(_06296_),
    .A3(_06321_),
    .A4(_06349_),
    .ZN(_06350_));
 NOR2_X2 _31447_ (.A1(_06350_),
    .A2(_05733_),
    .ZN(_06351_));
 AND4_X1 _31448_ (.A1(_05146_),
    .A2(_05438_),
    .A3(_05157_),
    .A4(_05227_),
    .ZN(_06352_));
 NOR2_X1 _31449_ (.A1(_05356_),
    .A2(_06352_),
    .ZN(_06353_));
 CLKBUF_X2 _31450_ (.A(_05338_),
    .Z(_06354_));
 NAND2_X1 _31451_ (.A1(_06354_),
    .A2(_05180_),
    .ZN(_06355_));
 AND3_X1 _31452_ (.A1(_05260_),
    .A2(_05327_),
    .A3(_05206_),
    .ZN(_06356_));
 AND2_X1 _31453_ (.A1(_05338_),
    .A2(_05176_),
    .ZN(_06357_));
 AOI211_X1 _31454_ (.A(_06356_),
    .B(_06357_),
    .C1(_05219_),
    .C2(_06354_),
    .ZN(_06359_));
 INV_X1 _31455_ (.A(_05238_),
    .ZN(_06360_));
 OAI21_X1 _31456_ (.A(_05347_),
    .B1(_06360_),
    .B2(_05306_),
    .ZN(_06361_));
 OAI21_X1 _31457_ (.A(_05347_),
    .B1(_05446_),
    .B2(_05359_),
    .ZN(_06362_));
 AND4_X1 _31458_ (.A1(_06355_),
    .A2(_06359_),
    .A3(_06361_),
    .A4(_06362_),
    .ZN(_06363_));
 OAI21_X1 _31459_ (.A(_05358_),
    .B1(_05430_),
    .B2(_05127_),
    .ZN(_06364_));
 AND2_X1 _31460_ (.A1(_05329_),
    .A2(_05462_),
    .ZN(_06365_));
 AND2_X1 _31461_ (.A1(_05329_),
    .A2(_05213_),
    .ZN(_06366_));
 AND2_X1 _31462_ (.A1(_05329_),
    .A2(_05252_),
    .ZN(_06367_));
 AND2_X1 _31463_ (.A1(_05328_),
    .A2(_05171_),
    .ZN(_06368_));
 NOR4_X1 _31464_ (.A1(_06365_),
    .A2(_06366_),
    .A3(_06367_),
    .A4(_06368_),
    .ZN(_06370_));
 AND4_X1 _31465_ (.A1(_06353_),
    .A2(_06363_),
    .A3(_06364_),
    .A4(_06370_),
    .ZN(_06371_));
 BUF_X2 _31466_ (.A(_05232_),
    .Z(_06372_));
 AND2_X1 _31467_ (.A1(_06372_),
    .A2(_05175_),
    .ZN(_06373_));
 INV_X1 _31468_ (.A(_05162_),
    .ZN(_06374_));
 OAI21_X1 _31469_ (.A(_05178_),
    .B1(_06374_),
    .B2(_05191_),
    .ZN(_06375_));
 AOI211_X1 _31470_ (.A(_06373_),
    .B(_06375_),
    .C1(_05171_),
    .C2(_05175_),
    .ZN(_06376_));
 INV_X1 _31471_ (.A(_05168_),
    .ZN(_06377_));
 AOI211_X1 _31472_ (.A(_06377_),
    .B(_05154_),
    .C1(_05164_),
    .C2(_05172_),
    .ZN(_06378_));
 INV_X1 _31473_ (.A(_05171_),
    .ZN(_06379_));
 AOI211_X1 _31474_ (.A(_06379_),
    .B(_05154_),
    .C1(_05164_),
    .C2(_05166_),
    .ZN(_06381_));
 NOR2_X1 _31475_ (.A1(_05154_),
    .A2(_05158_),
    .ZN(_06382_));
 NOR4_X1 _31476_ (.A1(_06378_),
    .A2(_06381_),
    .A3(_05480_),
    .A4(_06382_),
    .ZN(_06383_));
 BUF_X2 _31477_ (.A(_05187_),
    .Z(_06384_));
 AND2_X1 _31478_ (.A1(_06384_),
    .A2(_05284_),
    .ZN(_06385_));
 INV_X1 _31479_ (.A(_05235_),
    .ZN(_06386_));
 AOI21_X1 _31480_ (.A(_05195_),
    .B1(_05454_),
    .B2(_06386_),
    .ZN(_06387_));
 AND2_X1 _31481_ (.A1(_05150_),
    .A2(_05172_),
    .ZN(_06388_));
 AOI211_X1 _31482_ (.A(_06385_),
    .B(_06387_),
    .C1(_06388_),
    .C2(_06384_),
    .ZN(_06389_));
 INV_X1 _31483_ (.A(_05191_),
    .ZN(_06390_));
 OAI21_X1 _31484_ (.A(_05199_),
    .B1(_06390_),
    .B2(_05348_),
    .ZN(_06392_));
 AND4_X1 _31485_ (.A1(_06376_),
    .A2(_06383_),
    .A3(_06389_),
    .A4(_06392_),
    .ZN(_06393_));
 CLKBUF_X2 _31486_ (.A(_05286_),
    .Z(_06394_));
 AND3_X1 _31487_ (.A1(_06394_),
    .A2(_05168_),
    .A3(_05227_),
    .ZN(_06395_));
 AND3_X1 _31488_ (.A1(_05237_),
    .A2(_06394_),
    .A3(_05227_),
    .ZN(_06396_));
 AOI211_X1 _31489_ (.A(_06395_),
    .B(_06396_),
    .C1(_05235_),
    .C2(_05281_),
    .ZN(_06397_));
 NAND2_X1 _31490_ (.A1(_06390_),
    .A2(_05281_),
    .ZN(_06398_));
 OAI211_X1 _31491_ (.A(_06397_),
    .B(_06398_),
    .C1(_05294_),
    .C2(_05451_),
    .ZN(_06399_));
 OAI21_X1 _31492_ (.A(_05441_),
    .B1(_05389_),
    .B2(_05248_),
    .ZN(_06400_));
 OAI211_X1 _31493_ (.A(_06394_),
    .B(_05215_),
    .C1(_05127_),
    .C2(_05209_),
    .ZN(_06401_));
 NAND2_X1 _31494_ (.A1(_05441_),
    .A2(_05462_),
    .ZN(_06403_));
 NAND2_X1 _31495_ (.A1(_05441_),
    .A2(_05384_),
    .ZN(_06404_));
 NAND4_X1 _31496_ (.A1(_06400_),
    .A2(_06401_),
    .A3(_06403_),
    .A4(_06404_),
    .ZN(_06405_));
 OAI21_X1 _31497_ (.A(_05297_),
    .B1(_05235_),
    .B2(_06372_),
    .ZN(_06406_));
 OAI21_X1 _31498_ (.A(_05297_),
    .B1(_05261_),
    .B2(_05177_),
    .ZN(_06407_));
 INV_X1 _31499_ (.A(_06388_),
    .ZN(_06408_));
 OAI211_X1 _31500_ (.A(_06406_),
    .B(_06407_),
    .C1(_06408_),
    .C2(_05292_),
    .ZN(_06409_));
 BUF_X2 _31501_ (.A(_05150_),
    .Z(_06410_));
 NAND4_X1 _31502_ (.A1(_06394_),
    .A2(_06410_),
    .A3(_05138_),
    .A4(_05151_),
    .ZN(_06411_));
 NAND3_X1 _31503_ (.A1(_05311_),
    .A2(_05204_),
    .A3(_05190_),
    .ZN(_06412_));
 NAND4_X1 _31504_ (.A1(_05413_),
    .A2(_05392_),
    .A3(_06411_),
    .A4(_06412_),
    .ZN(_06414_));
 NOR4_X1 _31505_ (.A1(_06399_),
    .A2(_06405_),
    .A3(_06409_),
    .A4(_06414_),
    .ZN(_06415_));
 NAND2_X1 _31506_ (.A1(_05301_),
    .A2(_05220_),
    .ZN(_06416_));
 OAI211_X1 _31507_ (.A(_05221_),
    .B(_06416_),
    .C1(_05294_),
    .C2(_05239_),
    .ZN(_06417_));
 AOI21_X1 _31508_ (.A(_05239_),
    .B1(_05399_),
    .B2(_05436_),
    .ZN(_06418_));
 AND4_X1 _31509_ (.A1(_05215_),
    .A2(_05168_),
    .A3(_05146_),
    .A4(_05267_),
    .ZN(_06419_));
 NOR3_X1 _31510_ (.A1(_06417_),
    .A2(_06418_),
    .A3(_06419_),
    .ZN(_06420_));
 AND4_X1 _31511_ (.A1(_05124_),
    .A2(_05168_),
    .A3(_05151_),
    .A4(_05267_),
    .ZN(_06421_));
 AOI211_X1 _31512_ (.A(_05295_),
    .B(_05274_),
    .C1(_05164_),
    .C2(_05166_),
    .ZN(_06422_));
 AOI211_X1 _31513_ (.A(_06421_),
    .B(_06422_),
    .C1(_05332_),
    .C2(_05263_),
    .ZN(_06423_));
 OAI21_X1 _31514_ (.A(_05380_),
    .B1(_05250_),
    .B2(_05320_),
    .ZN(_06425_));
 NAND2_X1 _31515_ (.A1(_05316_),
    .A2(_05380_),
    .ZN(_06426_));
 NAND2_X1 _31516_ (.A1(_05209_),
    .A2(_05380_),
    .ZN(_06427_));
 AND4_X1 _31517_ (.A1(_05468_),
    .A2(_06425_),
    .A3(_06426_),
    .A4(_06427_),
    .ZN(_06428_));
 AND2_X1 _31518_ (.A1(_05458_),
    .A2(_05244_),
    .ZN(_06429_));
 AND2_X1 _31519_ (.A1(_05244_),
    .A2(_05462_),
    .ZN(_06430_));
 AND3_X1 _31520_ (.A1(_05384_),
    .A2(_05206_),
    .A3(_05267_),
    .ZN(_06431_));
 AND3_X1 _31521_ (.A1(_05446_),
    .A2(_05206_),
    .A3(_05267_),
    .ZN(_06432_));
 NOR4_X1 _31522_ (.A1(_06429_),
    .A2(_06430_),
    .A3(_06431_),
    .A4(_06432_),
    .ZN(_06433_));
 AND4_X1 _31523_ (.A1(_06420_),
    .A2(_06423_),
    .A3(_06428_),
    .A4(_06433_),
    .ZN(_06434_));
 NAND4_X1 _31524_ (.A1(_06371_),
    .A2(_06393_),
    .A3(_06415_),
    .A4(_06434_),
    .ZN(_06436_));
 NOR2_X2 _31525_ (.A1(_06436_),
    .A2(_05366_),
    .ZN(_06437_));
 XOR2_X2 _31526_ (.A(_06351_),
    .B(_06437_),
    .Z(_06438_));
 XNOR2_X1 _31527_ (.A(_05485_),
    .B(_06438_),
    .ZN(_06439_));
 NAND3_X1 _31528_ (.A1(_06170_),
    .A2(_06077_),
    .A3(_06037_),
    .ZN(_06440_));
 NAND3_X1 _31529_ (.A1(_06052_),
    .A2(_06077_),
    .A3(_06037_),
    .ZN(_06441_));
 NAND2_X1 _31530_ (.A1(_06440_),
    .A2(_06441_),
    .ZN(_06442_));
 INV_X1 _31531_ (.A(_06091_),
    .ZN(_06443_));
 AOI21_X1 _31532_ (.A(_06120_),
    .B1(_06098_),
    .B2(_06443_),
    .ZN(_06444_));
 AND2_X1 _31533_ (.A1(_06168_),
    .A2(_06119_),
    .ZN(_06445_));
 AOI211_X1 _31534_ (.A(_06442_),
    .B(_06444_),
    .C1(_06065_),
    .C2(_06445_),
    .ZN(_06447_));
 NAND2_X1 _31535_ (.A1(_06146_),
    .A2(_06078_),
    .ZN(_06448_));
 AND3_X1 _31536_ (.A1(_06078_),
    .A2(_06004_),
    .A3(_06027_),
    .ZN(_06449_));
 NOR2_X1 _31537_ (.A1(_06081_),
    .A2(_06449_),
    .ZN(_06450_));
 OAI21_X1 _31538_ (.A(_06078_),
    .B1(_06095_),
    .B2(_06048_),
    .ZN(_06451_));
 NAND4_X1 _31539_ (.A1(_06447_),
    .A2(_06448_),
    .A3(_06450_),
    .A4(_06451_),
    .ZN(_06452_));
 AND2_X1 _31540_ (.A1(_06048_),
    .A2(_06110_),
    .ZN(_06453_));
 INV_X1 _31541_ (.A(_06163_),
    .ZN(_06454_));
 INV_X1 _31542_ (.A(_06190_),
    .ZN(_06455_));
 NAND2_X1 _31543_ (.A1(_06454_),
    .A2(_06455_),
    .ZN(_06456_));
 INV_X1 _31544_ (.A(_06456_),
    .ZN(_06458_));
 INV_X1 _31545_ (.A(_06188_),
    .ZN(_06459_));
 AOI21_X1 _31546_ (.A(_06117_),
    .B1(_06458_),
    .B2(_06459_),
    .ZN(_06460_));
 AND2_X1 _31547_ (.A1(_06093_),
    .A2(_06110_),
    .ZN(_06461_));
 AND2_X1 _31548_ (.A1(_06052_),
    .A2(_06110_),
    .ZN(_06462_));
 OR4_X1 _31549_ (.A1(_06453_),
    .A2(_06460_),
    .A3(_06461_),
    .A4(_06462_),
    .ZN(_06463_));
 INV_X1 _31550_ (.A(_06090_),
    .ZN(_06464_));
 NAND2_X1 _31551_ (.A1(_05987_),
    .A2(_06005_),
    .ZN(_06465_));
 AND2_X1 _31552_ (.A1(_06043_),
    .A2(_16759_),
    .ZN(_06466_));
 INV_X1 _31553_ (.A(_06466_),
    .ZN(_06467_));
 AOI21_X1 _31554_ (.A(_06464_),
    .B1(_06465_),
    .B2(_06467_),
    .ZN(_06469_));
 AND2_X1 _31555_ (.A1(_06090_),
    .A2(_06170_),
    .ZN(_06470_));
 INV_X1 _31556_ (.A(_06470_),
    .ZN(_06471_));
 NAND3_X1 _31557_ (.A1(_06052_),
    .A2(_06172_),
    .A3(_06077_),
    .ZN(_06472_));
 OAI211_X1 _31558_ (.A(_06471_),
    .B(_06472_),
    .C1(_06464_),
    .C2(_06443_),
    .ZN(_06473_));
 NOR4_X1 _31559_ (.A1(_06452_),
    .A2(_06463_),
    .A3(_06469_),
    .A4(_06473_),
    .ZN(_06474_));
 NAND3_X1 _31560_ (.A1(_05996_),
    .A2(_06005_),
    .A3(_06198_),
    .ZN(_06475_));
 NAND3_X1 _31561_ (.A1(_05996_),
    .A2(_06005_),
    .A3(_05986_),
    .ZN(_06476_));
 NAND3_X1 _31562_ (.A1(_05996_),
    .A2(_06005_),
    .A3(_06032_),
    .ZN(_06477_));
 AND4_X1 _31563_ (.A1(_06001_),
    .A2(_06475_),
    .A3(_06476_),
    .A4(_06477_),
    .ZN(_06478_));
 AND2_X1 _31564_ (.A1(_06022_),
    .A2(_06085_),
    .ZN(_06480_));
 AND2_X1 _31565_ (.A1(_06012_),
    .A2(_16760_),
    .ZN(_06481_));
 CLKBUF_X2 _31566_ (.A(_06481_),
    .Z(_06482_));
 AND2_X1 _31567_ (.A1(_06022_),
    .A2(_06482_),
    .ZN(_06483_));
 AND2_X1 _31568_ (.A1(_06004_),
    .A2(_06045_),
    .ZN(_06484_));
 AND2_X1 _31569_ (.A1(_06022_),
    .A2(_06484_),
    .ZN(_06485_));
 AND2_X1 _31570_ (.A1(_06022_),
    .A2(_06143_),
    .ZN(_06486_));
 NOR4_X1 _31571_ (.A1(_06480_),
    .A2(_06483_),
    .A3(_06485_),
    .A4(_06486_),
    .ZN(_06487_));
 AND3_X1 _31572_ (.A1(_05996_),
    .A2(_06032_),
    .A3(_06013_),
    .ZN(_06488_));
 AND2_X1 _31573_ (.A1(_06095_),
    .A2(_05996_),
    .ZN(_06489_));
 AND2_X1 _31574_ (.A1(_06211_),
    .A2(_05996_),
    .ZN(_06491_));
 AND2_X1 _31575_ (.A1(_06048_),
    .A2(_05996_),
    .ZN(_06492_));
 NOR4_X1 _31576_ (.A1(_06488_),
    .A2(_06489_),
    .A3(_06491_),
    .A4(_06492_),
    .ZN(_06493_));
 OAI21_X1 _31577_ (.A(_06038_),
    .B1(_06019_),
    .B2(_06124_),
    .ZN(_06494_));
 INV_X1 _31578_ (.A(_06067_),
    .ZN(_06495_));
 OAI21_X1 _31579_ (.A(_06063_),
    .B1(_06495_),
    .B2(_06188_),
    .ZN(_06496_));
 OAI211_X1 _31580_ (.A(_06063_),
    .B(_06013_),
    .C1(_06044_),
    .C2(_06009_),
    .ZN(_06497_));
 OAI211_X1 _31581_ (.A(_06063_),
    .B(_06058_),
    .C1(_06044_),
    .C2(_06045_),
    .ZN(_06498_));
 AND4_X1 _31582_ (.A1(_06494_),
    .A2(_06496_),
    .A3(_06497_),
    .A4(_06498_),
    .ZN(_06499_));
 AND4_X1 _31583_ (.A1(_06478_),
    .A2(_06487_),
    .A3(_06493_),
    .A4(_06499_),
    .ZN(_06500_));
 OAI21_X1 _31584_ (.A(_06136_),
    .B1(_06019_),
    .B2(_06466_),
    .ZN(_06502_));
 OAI21_X1 _31585_ (.A(_06136_),
    .B1(_06099_),
    .B2(_06482_),
    .ZN(_06503_));
 OAI21_X1 _31586_ (.A(_06136_),
    .B1(_06106_),
    .B2(_06085_),
    .ZN(_06504_));
 AND3_X1 _31587_ (.A1(_06502_),
    .A2(_06503_),
    .A3(_06504_),
    .ZN(_06505_));
 INV_X1 _31588_ (.A(_06151_),
    .ZN(_06506_));
 AOI21_X1 _31589_ (.A(_06174_),
    .B1(_06455_),
    .B2(_06506_),
    .ZN(_06507_));
 AOI21_X1 _31590_ (.A(_06174_),
    .B1(_06098_),
    .B2(_06443_),
    .ZN(_06508_));
 NAND2_X1 _31591_ (.A1(_06125_),
    .A2(_06058_),
    .ZN(_06509_));
 NOR2_X1 _31592_ (.A1(_06509_),
    .A2(_06198_),
    .ZN(_06510_));
 AOI211_X1 _31593_ (.A(_06507_),
    .B(_06508_),
    .C1(_06166_),
    .C2(_06510_),
    .ZN(_06511_));
 AND2_X1 _31594_ (.A1(_06495_),
    .A2(_06145_),
    .ZN(_06513_));
 INV_X1 _31595_ (.A(_06481_),
    .ZN(_06514_));
 OAI21_X1 _31596_ (.A(_06157_),
    .B1(_06161_),
    .B2(_06514_),
    .ZN(_06515_));
 AOI211_X1 _31597_ (.A(_06513_),
    .B(_06515_),
    .C1(_06484_),
    .C2(_06145_),
    .ZN(_06516_));
 AND2_X1 _31598_ (.A1(_05990_),
    .A2(_06179_),
    .ZN(_06517_));
 NAND2_X1 _31599_ (.A1(_06179_),
    .A2(_06466_),
    .ZN(_06518_));
 NAND4_X1 _31600_ (.A1(_06158_),
    .A2(_06005_),
    .A3(_05986_),
    .A4(_06183_),
    .ZN(_06519_));
 NAND2_X1 _31601_ (.A1(_06518_),
    .A2(_06519_),
    .ZN(_06520_));
 NOR3_X2 _31602_ (.A1(_06150_),
    .A2(_16761_),
    .A3(_06011_),
    .ZN(_06521_));
 AND2_X1 _31603_ (.A1(_06521_),
    .A2(_05987_),
    .ZN(_06522_));
 AOI211_X1 _31604_ (.A(_06517_),
    .B(_06520_),
    .C1(_06180_),
    .C2(_06522_),
    .ZN(_06524_));
 AND4_X1 _31605_ (.A1(_06505_),
    .A2(_06511_),
    .A3(_06516_),
    .A4(_06524_),
    .ZN(_06525_));
 OAI211_X1 _31606_ (.A(_06202_),
    .B(_06058_),
    .C1(_06198_),
    .C2(_06032_),
    .ZN(_06526_));
 OAI21_X1 _31607_ (.A(_06202_),
    .B1(_06146_),
    .B2(_06223_),
    .ZN(_06527_));
 NAND4_X1 _31608_ (.A1(_06013_),
    .A2(_06195_),
    .A3(_06009_),
    .A4(_06183_),
    .ZN(_06528_));
 AND3_X1 _31609_ (.A1(_06526_),
    .A2(_06527_),
    .A3(_06528_),
    .ZN(_06529_));
 NAND2_X1 _31610_ (.A1(_06101_),
    .A2(_06209_),
    .ZN(_06530_));
 AND2_X1 _31611_ (.A1(_06099_),
    .A2(_06208_),
    .ZN(_06531_));
 AND2_X1 _31612_ (.A1(_06209_),
    .A2(_06093_),
    .ZN(_06532_));
 NOR2_X1 _31613_ (.A1(_06531_),
    .A2(_06532_),
    .ZN(_06533_));
 NAND2_X1 _31614_ (.A1(_06209_),
    .A2(_06075_),
    .ZN(_06535_));
 AND2_X1 _31615_ (.A1(_06209_),
    .A2(_06000_),
    .ZN(_06536_));
 INV_X1 _31616_ (.A(_06536_),
    .ZN(_06537_));
 AND4_X1 _31617_ (.A1(_06530_),
    .A2(_06533_),
    .A3(_06535_),
    .A4(_06537_),
    .ZN(_06538_));
 INV_X1 _31618_ (.A(_06221_),
    .ZN(_06539_));
 INV_X1 _31619_ (.A(_06102_),
    .ZN(_06540_));
 AOI21_X1 _31620_ (.A(_06539_),
    .B1(_06459_),
    .B2(_06540_),
    .ZN(_06541_));
 AND3_X1 _31621_ (.A1(_06221_),
    .A2(_05987_),
    .A3(_06521_),
    .ZN(_06542_));
 AND2_X1 _31622_ (.A1(_06221_),
    .A2(_06170_),
    .ZN(_06543_));
 NOR4_X1 _31623_ (.A1(_06541_),
    .A2(_06542_),
    .A3(_06222_),
    .A4(_06543_),
    .ZN(_06544_));
 NAND2_X1 _31624_ (.A1(_06196_),
    .A2(_06103_),
    .ZN(_06546_));
 OAI21_X1 _31625_ (.A(_06196_),
    .B1(_06048_),
    .B2(_06211_),
    .ZN(_06547_));
 NAND2_X1 _31626_ (.A1(_06196_),
    .A2(_06128_),
    .ZN(_06548_));
 NAND2_X1 _31627_ (.A1(_06196_),
    .A2(_06099_),
    .ZN(_06549_));
 AND4_X1 _31628_ (.A1(_06546_),
    .A2(_06547_),
    .A3(_06548_),
    .A4(_06549_),
    .ZN(_06550_));
 AND4_X1 _31629_ (.A1(_06529_),
    .A2(_06538_),
    .A3(_06544_),
    .A4(_06550_),
    .ZN(_06551_));
 NAND4_X1 _31630_ (.A1(_06474_),
    .A2(_06500_),
    .A3(_06525_),
    .A4(_06551_),
    .ZN(_06552_));
 NOR2_X2 _31631_ (.A1(_06552_),
    .A2(_06232_),
    .ZN(_06553_));
 XNOR2_X1 _31632_ (.A(_06553_),
    .B(_00989_),
    .ZN(_06554_));
 AND3_X1 _31633_ (.A1(_05908_),
    .A2(_05778_),
    .A3(_05743_),
    .ZN(_06555_));
 AOI21_X1 _31634_ (.A(_06555_),
    .B1(_05969_),
    .B2(_05939_),
    .ZN(_06557_));
 AND3_X1 _31635_ (.A1(_05938_),
    .A2(_05743_),
    .A3(_05759_),
    .ZN(_06558_));
 BUF_X2 _31636_ (.A(_05917_),
    .Z(_06559_));
 AOI21_X1 _31637_ (.A(_06558_),
    .B1(_06559_),
    .B2(_05967_),
    .ZN(_06560_));
 BUF_X2 _31638_ (.A(_05870_),
    .Z(_06561_));
 AOI22_X1 _31639_ (.A1(_05857_),
    .A2(_05883_),
    .B1(_06561_),
    .B2(_06559_),
    .ZN(_06562_));
 AOI22_X1 _31640_ (.A1(_05864_),
    .A2(_05909_),
    .B1(_05783_),
    .B2(_05883_),
    .ZN(_06563_));
 AND4_X1 _31641_ (.A1(_06557_),
    .A2(_06560_),
    .A3(_06562_),
    .A4(_06563_),
    .ZN(_06564_));
 AND2_X1 _31642_ (.A1(_05972_),
    .A2(_05765_),
    .ZN(_06565_));
 INV_X1 _31643_ (.A(_05771_),
    .ZN(_06566_));
 AND2_X1 _31644_ (.A1(_05787_),
    .A2(_05763_),
    .ZN(_06568_));
 INV_X1 _31645_ (.A(_06568_),
    .ZN(_06569_));
 AND2_X1 _31646_ (.A1(_05759_),
    .A2(_05745_),
    .ZN(_06570_));
 NAND3_X1 _31647_ (.A1(_06570_),
    .A2(_05849_),
    .A3(_05802_),
    .ZN(_06571_));
 BUF_X2 _31648_ (.A(_16800_),
    .Z(_06572_));
 OAI22_X1 _31649_ (.A1(_06566_),
    .A2(_06569_),
    .B1(_06571_),
    .B2(_06572_),
    .ZN(_06573_));
 AOI211_X1 _31650_ (.A(_06565_),
    .B(_06573_),
    .C1(_05931_),
    .C2(_05774_),
    .ZN(_06574_));
 AND2_X2 _31651_ (.A1(_05821_),
    .A2(_05759_),
    .ZN(_06575_));
 NAND3_X1 _31652_ (.A1(_05952_),
    .A2(_06575_),
    .A3(_05872_),
    .ZN(_06576_));
 OAI21_X1 _31653_ (.A(_05765_),
    .B1(_05860_),
    .B2(_05909_),
    .ZN(_06577_));
 AND2_X1 _31654_ (.A1(_06576_),
    .A2(_06577_),
    .ZN(_06579_));
 OAI21_X1 _31655_ (.A(_05785_),
    .B1(_05821_),
    .B2(_16801_),
    .ZN(_06580_));
 AND3_X1 _31656_ (.A1(_05748_),
    .A2(_05749_),
    .A3(_05785_),
    .ZN(_06581_));
 AOI21_X1 _31657_ (.A(_16802_),
    .B1(_05780_),
    .B2(_05737_),
    .ZN(_06582_));
 AOI22_X1 _31658_ (.A1(_06580_),
    .A2(_06581_),
    .B1(_05828_),
    .B2(_06582_),
    .ZN(_06583_));
 AND4_X1 _31659_ (.A1(_06564_),
    .A2(_06574_),
    .A3(_06579_),
    .A4(_06583_),
    .ZN(_06584_));
 NOR2_X1 _31660_ (.A1(_05916_),
    .A2(_05880_),
    .ZN(_06585_));
 AND2_X1 _31661_ (.A1(_05744_),
    .A2(_05967_),
    .ZN(_06586_));
 AND2_X1 _31662_ (.A1(_05827_),
    .A2(_05969_),
    .ZN(_06587_));
 AND2_X1 _31663_ (.A1(_06568_),
    .A2(_05883_),
    .ZN(_06588_));
 NOR4_X1 _31664_ (.A1(_05875_),
    .A2(_06586_),
    .A3(_06587_),
    .A4(_06588_),
    .ZN(_06590_));
 INV_X1 _31665_ (.A(_05967_),
    .ZN(_06591_));
 NAND2_X1 _31666_ (.A1(_05747_),
    .A2(_05851_),
    .ZN(_06592_));
 NOR2_X1 _31667_ (.A1(_06591_),
    .A2(_06592_),
    .ZN(_06593_));
 INV_X1 _31668_ (.A(_06593_),
    .ZN(_06594_));
 AND2_X1 _31669_ (.A1(_05787_),
    .A2(_16799_),
    .ZN(_06595_));
 AOI22_X1 _31670_ (.A1(_05886_),
    .A2(_06575_),
    .B1(_06595_),
    .B2(_05939_),
    .ZN(_06596_));
 AND4_X1 _31671_ (.A1(_06585_),
    .A2(_06590_),
    .A3(_06594_),
    .A4(_06596_),
    .ZN(_06597_));
 INV_X1 _31672_ (.A(_05899_),
    .ZN(_06598_));
 INV_X1 _31673_ (.A(_05963_),
    .ZN(_06599_));
 INV_X1 _31674_ (.A(_05867_),
    .ZN(_06601_));
 AOI21_X1 _31675_ (.A(_06598_),
    .B1(_06599_),
    .B2(_06601_),
    .ZN(_06602_));
 INV_X1 _31676_ (.A(_06602_),
    .ZN(_06603_));
 BUF_X2 _31677_ (.A(_05925_),
    .Z(_06604_));
 NOR2_X2 _31678_ (.A1(_05822_),
    .A2(_05767_),
    .ZN(_06605_));
 OAI21_X1 _31679_ (.A(_06604_),
    .B1(_06605_),
    .B2(_05855_),
    .ZN(_06606_));
 NAND2_X1 _31680_ (.A1(_05872_),
    .A2(_05739_),
    .ZN(_06607_));
 NOR2_X1 _31681_ (.A1(_06607_),
    .A2(_05763_),
    .ZN(_06608_));
 CLKBUF_X2 _31682_ (.A(_05837_),
    .Z(_06609_));
 OAI21_X1 _31683_ (.A(_06561_),
    .B1(_06608_),
    .B2(_06609_),
    .ZN(_06610_));
 OAI21_X1 _31684_ (.A(_05972_),
    .B1(_05834_),
    .B2(_05794_),
    .ZN(_06612_));
 NAND3_X1 _31685_ (.A1(_05972_),
    .A2(_05850_),
    .A3(_06609_),
    .ZN(_06613_));
 NAND2_X1 _31686_ (.A1(_05823_),
    .A2(_05958_),
    .ZN(_06614_));
 AND3_X1 _31687_ (.A1(_06612_),
    .A2(_06613_),
    .A3(_06614_),
    .ZN(_06615_));
 AND4_X1 _31688_ (.A1(_06603_),
    .A2(_06606_),
    .A3(_06610_),
    .A4(_06615_),
    .ZN(_06616_));
 AND2_X1 _31689_ (.A1(_05925_),
    .A2(_05866_),
    .ZN(_06617_));
 AND2_X1 _31690_ (.A1(_05739_),
    .A2(_16799_),
    .ZN(_06618_));
 AND2_X1 _31691_ (.A1(_06618_),
    .A2(_05803_),
    .ZN(_06619_));
 AND3_X1 _31692_ (.A1(_05831_),
    .A2(_05756_),
    .A3(_05749_),
    .ZN(_06620_));
 NOR4_X1 _31693_ (.A1(_06617_),
    .A2(_06619_),
    .A3(_05805_),
    .A4(_06620_),
    .ZN(_06621_));
 AND2_X1 _31694_ (.A1(_05843_),
    .A2(_05876_),
    .ZN(_06623_));
 AND2_X1 _31695_ (.A1(_05952_),
    .A2(_05837_),
    .ZN(_06624_));
 AND2_X1 _31696_ (.A1(_05866_),
    .A2(_05750_),
    .ZN(_06625_));
 AND3_X1 _31697_ (.A1(_05829_),
    .A2(_05849_),
    .A3(_05748_),
    .ZN(_06626_));
 NOR4_X1 _31698_ (.A1(_06623_),
    .A2(_06624_),
    .A3(_06625_),
    .A4(_06626_),
    .ZN(_06627_));
 AND2_X1 _31699_ (.A1(_05811_),
    .A2(_05900_),
    .ZN(_06628_));
 AND2_X1 _31700_ (.A1(_05794_),
    .A2(_05938_),
    .ZN(_06629_));
 NOR3_X1 _31701_ (.A1(_05927_),
    .A2(_06628_),
    .A3(_06629_),
    .ZN(_06630_));
 AND2_X1 _31702_ (.A1(_05925_),
    .A2(_05789_),
    .ZN(_06631_));
 AND2_X1 _31703_ (.A1(_05789_),
    .A2(_05909_),
    .ZN(_06632_));
 AND2_X1 _31704_ (.A1(_05794_),
    .A2(_05883_),
    .ZN(_06634_));
 AND2_X1 _31705_ (.A1(_05909_),
    .A2(_05791_),
    .ZN(_06635_));
 NOR4_X1 _31706_ (.A1(_06631_),
    .A2(_06632_),
    .A3(_06634_),
    .A4(_06635_),
    .ZN(_06636_));
 AND4_X1 _31707_ (.A1(_06621_),
    .A2(_06627_),
    .A3(_06630_),
    .A4(_06636_),
    .ZN(_06637_));
 NAND4_X1 _31708_ (.A1(_06584_),
    .A2(_06597_),
    .A3(_06616_),
    .A4(_06637_),
    .ZN(_06638_));
 NOR3_X1 _31709_ (.A1(_05744_),
    .A2(_06595_),
    .A3(_06570_),
    .ZN(_06639_));
 INV_X1 _31710_ (.A(_05957_),
    .ZN(_06640_));
 NOR2_X1 _31711_ (.A1(_06639_),
    .A2(_06640_),
    .ZN(_06641_));
 NAND4_X1 _31712_ (.A1(_05848_),
    .A2(_05977_),
    .A3(_05849_),
    .A4(_05850_),
    .ZN(_06642_));
 INV_X1 _31713_ (.A(_05842_),
    .ZN(_06643_));
 OAI21_X1 _31714_ (.A(_06642_),
    .B1(_06643_),
    .B2(_05953_),
    .ZN(_06645_));
 INV_X1 _31715_ (.A(_05751_),
    .ZN(_06646_));
 INV_X1 _31716_ (.A(_05855_),
    .ZN(_06647_));
 AOI22_X1 _31717_ (.A1(_05977_),
    .A2(_05746_),
    .B1(_06572_),
    .B2(_05785_),
    .ZN(_06648_));
 AOI21_X1 _31718_ (.A(_06646_),
    .B1(_06647_),
    .B2(_06648_),
    .ZN(_06649_));
 NOR3_X1 _31719_ (.A1(_06646_),
    .A2(_05767_),
    .A3(_05822_),
    .ZN(_06650_));
 NOR4_X1 _31720_ (.A1(_06641_),
    .A2(_06645_),
    .A3(_06649_),
    .A4(_06650_),
    .ZN(_06651_));
 NAND3_X1 _31721_ (.A1(_05823_),
    .A2(_05872_),
    .A3(_05809_),
    .ZN(_06652_));
 NAND2_X1 _31722_ (.A1(_05931_),
    .A2(_05809_),
    .ZN(_06653_));
 NAND2_X1 _31723_ (.A1(_06652_),
    .A2(_06653_),
    .ZN(_06654_));
 INV_X1 _31724_ (.A(_06654_),
    .ZN(_06656_));
 OAI21_X1 _31725_ (.A(_05774_),
    .B1(_05855_),
    .B2(_05857_),
    .ZN(_06657_));
 NAND4_X1 _31726_ (.A1(_05977_),
    .A2(_05849_),
    .A3(_05850_),
    .A4(_05748_),
    .ZN(_06658_));
 OAI21_X1 _31727_ (.A(_05861_),
    .B1(_05969_),
    .B2(_05794_),
    .ZN(_06659_));
 NOR3_X1 _31728_ (.A1(_05743_),
    .A2(_05785_),
    .A3(_16801_),
    .ZN(_06660_));
 NAND2_X1 _31729_ (.A1(_06660_),
    .A2(_05828_),
    .ZN(_06661_));
 INV_X1 _31730_ (.A(_05887_),
    .ZN(_06662_));
 NAND4_X1 _31731_ (.A1(_06662_),
    .A2(_05848_),
    .A3(_05851_),
    .A4(_05849_),
    .ZN(_06663_));
 AND4_X1 _31732_ (.A1(_06658_),
    .A2(_06659_),
    .A3(_06661_),
    .A4(_06663_),
    .ZN(_06664_));
 NAND4_X1 _31733_ (.A1(_06651_),
    .A2(_06656_),
    .A3(_06657_),
    .A4(_06664_),
    .ZN(_06665_));
 NOR2_X2 _31734_ (.A1(_06638_),
    .A2(_06665_),
    .ZN(_06667_));
 INV_X1 _31735_ (.A(_06667_),
    .ZN(_06668_));
 XNOR2_X2 _31736_ (.A(_06668_),
    .B(_05983_),
    .ZN(_06669_));
 XOR2_X1 _31737_ (.A(_06554_),
    .B(_06669_),
    .Z(_06670_));
 XNOR2_X1 _31738_ (.A(_06439_),
    .B(_06670_),
    .ZN(_06671_));
 MUX2_X1 _31739_ (.A(_06239_),
    .B(_06671_),
    .S(_05069_),
    .Z(_00701_));
 MUX2_X1 _31740_ (.A(_16942_),
    .B(_16814_),
    .S(_06237_),
    .Z(_00739_));
 MUX2_X1 _31741_ (.A(_16943_),
    .B(_16815_),
    .S(_06237_),
    .Z(_00740_));
 MUX2_X1 _31742_ (.A(_16944_),
    .B(_16816_),
    .S(_06237_),
    .Z(_00741_));
 MUX2_X1 _31743_ (.A(_16945_),
    .B(_16817_),
    .S(_06237_),
    .Z(_00742_));
 MUX2_X1 _31744_ (.A(_16947_),
    .B(_16819_),
    .S(_06237_),
    .Z(_00744_));
 BUF_X2 _31745_ (.A(_05104_),
    .Z(_06673_));
 MUX2_X1 _31746_ (.A(_16948_),
    .B(_16820_),
    .S(_06673_),
    .Z(_00745_));
 MUX2_X1 _31747_ (.A(_16949_),
    .B(_16821_),
    .S(_06673_),
    .Z(_00746_));
 MUX2_X1 _31748_ (.A(_16950_),
    .B(_16822_),
    .S(_06673_),
    .Z(_00747_));
 MUX2_X1 _31749_ (.A(_16951_),
    .B(_16823_),
    .S(_06673_),
    .Z(_00748_));
 MUX2_X1 _31750_ (.A(_16952_),
    .B(_16824_),
    .S(_06673_),
    .Z(_00749_));
 XOR2_X1 _31751_ (.A(_17121_),
    .B(_17060_),
    .Z(_06674_));
 INV_X1 _31752_ (.A(_05689_),
    .ZN(_06675_));
 AOI21_X1 _31753_ (.A(_05663_),
    .B1(_05565_),
    .B2(_06675_),
    .ZN(_06676_));
 AOI21_X1 _31754_ (.A(_05663_),
    .B1(_06341_),
    .B2(_06249_),
    .ZN(_06678_));
 AND4_X1 _31755_ (.A1(_05593_),
    .A2(_05638_),
    .A3(_05589_),
    .A4(_06309_),
    .ZN(_06679_));
 OR4_X1 _31756_ (.A1(_05668_),
    .A2(_06676_),
    .A3(_06678_),
    .A4(_06679_),
    .ZN(_06680_));
 OAI211_X1 _31757_ (.A(_05651_),
    .B(_16722_),
    .C1(_05711_),
    .C2(_05518_),
    .ZN(_06681_));
 OAI21_X1 _31758_ (.A(_05651_),
    .B1(_05690_),
    .B2(_05521_),
    .ZN(_06682_));
 OAI21_X1 _31759_ (.A(_05651_),
    .B1(_05619_),
    .B2(_05616_),
    .ZN(_06683_));
 NAND3_X1 _31760_ (.A1(_06681_),
    .A2(_06682_),
    .A3(_06683_),
    .ZN(_06684_));
 OAI211_X1 _31761_ (.A(_06272_),
    .B(_06312_),
    .C1(_05633_),
    .C2(_05705_),
    .ZN(_06685_));
 NAND3_X1 _31762_ (.A1(_05575_),
    .A2(_06272_),
    .A3(_06312_),
    .ZN(_06686_));
 OAI211_X1 _31763_ (.A(_06685_),
    .B(_06686_),
    .C1(_06261_),
    .C2(_05649_),
    .ZN(_06687_));
 AND2_X1 _31764_ (.A1(_05672_),
    .A2(_06275_),
    .ZN(_06689_));
 INV_X1 _31765_ (.A(_06689_),
    .ZN(_06690_));
 OAI21_X1 _31766_ (.A(_05673_),
    .B1(_05699_),
    .B2(_05521_),
    .ZN(_06691_));
 NOR2_X1 _31767_ (.A1(_05605_),
    .A2(_05701_),
    .ZN(_06692_));
 OAI211_X1 _31768_ (.A(_06690_),
    .B(_06691_),
    .C1(_06692_),
    .C2(_06319_),
    .ZN(_06693_));
 NOR4_X1 _31769_ (.A1(_06680_),
    .A2(_06684_),
    .A3(_06687_),
    .A4(_06693_),
    .ZN(_06694_));
 AND3_X1 _31770_ (.A1(_05557_),
    .A2(_06272_),
    .A3(_05714_),
    .ZN(_06695_));
 AND2_X1 _31771_ (.A1(_05696_),
    .A2(_06346_),
    .ZN(_06696_));
 NOR2_X1 _31772_ (.A1(_06302_),
    .A2(_05535_),
    .ZN(_06697_));
 AOI211_X1 _31773_ (.A(_06695_),
    .B(_06696_),
    .C1(_05696_),
    .C2(_06697_),
    .ZN(_06698_));
 OAI21_X1 _31774_ (.A(_05696_),
    .B1(_05646_),
    .B2(_05543_),
    .ZN(_06700_));
 AND3_X1 _31775_ (.A1(_06698_),
    .A2(_06323_),
    .A3(_06700_),
    .ZN(_06701_));
 NAND2_X1 _31776_ (.A1(_06271_),
    .A2(_06343_),
    .ZN(_06702_));
 INV_X1 _31777_ (.A(_05618_),
    .ZN(_06703_));
 INV_X1 _31778_ (.A(_06268_),
    .ZN(_06704_));
 NAND2_X1 _31779_ (.A1(_06703_),
    .A2(_06704_),
    .ZN(_06705_));
 OAI21_X1 _31780_ (.A(_05722_),
    .B1(_06705_),
    .B2(_05690_),
    .ZN(_06706_));
 OAI21_X1 _31781_ (.A(_06343_),
    .B1(_06697_),
    .B2(_05521_),
    .ZN(_06707_));
 OAI21_X1 _31782_ (.A(_05722_),
    .B1(_05703_),
    .B2(_05692_),
    .ZN(_06708_));
 AND4_X1 _31783_ (.A1(_06702_),
    .A2(_06706_),
    .A3(_06707_),
    .A4(_06708_),
    .ZN(_06709_));
 BUF_X2 _31784_ (.A(_05710_),
    .Z(_06711_));
 AND2_X1 _31785_ (.A1(_06711_),
    .A2(_05543_),
    .ZN(_06712_));
 INV_X1 _31786_ (.A(_05520_),
    .ZN(_06713_));
 AOI21_X1 _31787_ (.A(_05718_),
    .B1(_06675_),
    .B2(_06713_),
    .ZN(_06714_));
 OAI22_X1 _31788_ (.A1(_05711_),
    .A2(_05592_),
    .B1(_05666_),
    .B2(_05502_),
    .ZN(_06715_));
 AOI211_X1 _31789_ (.A(_06712_),
    .B(_06714_),
    .C1(_06711_),
    .C2(_06715_),
    .ZN(_06716_));
 NAND4_X1 _31790_ (.A1(_06694_),
    .A2(_06701_),
    .A3(_06709_),
    .A4(_06716_),
    .ZN(_06717_));
 NAND2_X1 _31791_ (.A1(_05626_),
    .A2(_05619_),
    .ZN(_06718_));
 AOI211_X1 _31792_ (.A(_06263_),
    .B(_05598_),
    .C1(_05657_),
    .C2(_05666_),
    .ZN(_06719_));
 AND2_X1 _31793_ (.A1(_05606_),
    .A2(_05646_),
    .ZN(_06720_));
 AND4_X1 _31794_ (.A1(_06285_),
    .A2(_05606_),
    .A3(_05657_),
    .A4(_05666_),
    .ZN(_06722_));
 NAND2_X1 _31795_ (.A1(_05699_),
    .A2(_05606_),
    .ZN(_06723_));
 NAND2_X1 _31796_ (.A1(_05597_),
    .A2(_06267_),
    .ZN(_06724_));
 NAND2_X1 _31797_ (.A1(_06723_),
    .A2(_06724_),
    .ZN(_06725_));
 NOR4_X1 _31798_ (.A1(_06719_),
    .A2(_06720_),
    .A3(_06722_),
    .A4(_06725_),
    .ZN(_06726_));
 OAI21_X1 _31799_ (.A(_05626_),
    .B1(_05701_),
    .B2(_05705_),
    .ZN(_06727_));
 AND4_X1 _31800_ (.A1(_06718_),
    .A2(_06726_),
    .A3(_05627_),
    .A4(_06727_),
    .ZN(_06728_));
 AND2_X1 _31801_ (.A1(_05536_),
    .A2(_05504_),
    .ZN(_06729_));
 OAI21_X1 _31802_ (.A(_05554_),
    .B1(_06729_),
    .B2(_05570_),
    .ZN(_06730_));
 AND2_X1 _31803_ (.A1(_05505_),
    .A2(_05572_),
    .ZN(_06731_));
 OAI21_X1 _31804_ (.A(_06251_),
    .B1(_06731_),
    .B2(_05692_),
    .ZN(_06733_));
 NAND4_X1 _31805_ (.A1(_06309_),
    .A2(_05715_),
    .A3(_05506_),
    .A4(_05711_),
    .ZN(_06734_));
 NAND4_X1 _31806_ (.A1(_06251_),
    .A2(_06291_),
    .A3(_05537_),
    .A4(_05532_),
    .ZN(_06735_));
 AND3_X1 _31807_ (.A1(_06733_),
    .A2(_06734_),
    .A3(_06735_),
    .ZN(_06736_));
 NAND2_X1 _31808_ (.A1(_05554_),
    .A2(_05686_),
    .ZN(_06737_));
 OAI21_X1 _31809_ (.A(_05554_),
    .B1(_05690_),
    .B2(_05521_),
    .ZN(_06738_));
 AND4_X1 _31810_ (.A1(_06730_),
    .A2(_06736_),
    .A3(_06737_),
    .A4(_06738_),
    .ZN(_06739_));
 OAI21_X1 _31811_ (.A(_05583_),
    .B1(_05699_),
    .B2(_05644_),
    .ZN(_06740_));
 OAI21_X1 _31812_ (.A(_06266_),
    .B1(_05699_),
    .B2(_05619_),
    .ZN(_06741_));
 OAI21_X1 _31813_ (.A(_06266_),
    .B1(_06275_),
    .B2(_05692_),
    .ZN(_06742_));
 OAI21_X1 _31814_ (.A(_05583_),
    .B1(_06275_),
    .B2(_06346_),
    .ZN(_06744_));
 AND4_X1 _31815_ (.A1(_06740_),
    .A2(_06741_),
    .A3(_06742_),
    .A4(_06744_),
    .ZN(_06745_));
 OAI21_X1 _31816_ (.A(_05541_),
    .B1(_05564_),
    .B2(_05619_),
    .ZN(_06746_));
 OAI21_X1 _31817_ (.A(_05541_),
    .B1(_05633_),
    .B2(_05705_),
    .ZN(_06747_));
 NAND3_X1 _31818_ (.A1(_05575_),
    .A2(_06272_),
    .A3(_05506_),
    .ZN(_06748_));
 NAND3_X1 _31819_ (.A1(_06746_),
    .A2(_06747_),
    .A3(_06748_),
    .ZN(_06749_));
 OAI21_X1 _31820_ (.A(_05490_),
    .B1(_05570_),
    .B2(_05575_),
    .ZN(_06750_));
 NAND3_X1 _31821_ (.A1(_05491_),
    .A2(_06285_),
    .A3(_05713_),
    .ZN(_06751_));
 NAND2_X1 _31822_ (.A1(_06750_),
    .A2(_06751_),
    .ZN(_06752_));
 NOR3_X1 _31823_ (.A1(_05510_),
    .A2(_05535_),
    .A3(_05568_),
    .ZN(_06753_));
 NOR4_X1 _31824_ (.A1(_06749_),
    .A2(_06752_),
    .A3(_06753_),
    .A4(_05523_),
    .ZN(_06755_));
 NAND4_X1 _31825_ (.A1(_06728_),
    .A2(_06739_),
    .A3(_06745_),
    .A4(_06755_),
    .ZN(_06756_));
 NOR2_X2 _31826_ (.A1(_06717_),
    .A2(_06756_),
    .ZN(_06757_));
 OAI21_X1 _31827_ (.A(_05244_),
    .B1(_05430_),
    .B2(_05301_),
    .ZN(_06758_));
 NOR2_X1 _31828_ (.A1(_05256_),
    .A2(_05141_),
    .ZN(_06759_));
 OR2_X1 _31829_ (.A1(_05255_),
    .A2(_06759_),
    .ZN(_06760_));
 OAI21_X1 _31830_ (.A(_05263_),
    .B1(_06372_),
    .B2(_05256_),
    .ZN(_06761_));
 OAI21_X1 _31831_ (.A(_05263_),
    .B1(_05250_),
    .B2(_05252_),
    .ZN(_06762_));
 AND4_X1 _31832_ (.A1(_06758_),
    .A2(_06760_),
    .A3(_06761_),
    .A4(_06762_),
    .ZN(_06763_));
 AND2_X1 _31833_ (.A1(_06354_),
    .A2(_05384_),
    .ZN(_06764_));
 AOI21_X1 _31834_ (.A(_06764_),
    .B1(_06360_),
    .B2(_06354_),
    .ZN(_06766_));
 BUF_X2 _31835_ (.A(_05206_),
    .Z(_06767_));
 NAND3_X1 _31836_ (.A1(_05219_),
    .A2(_05438_),
    .A3(_06767_),
    .ZN(_06768_));
 OAI211_X1 _31837_ (.A(_06766_),
    .B(_06768_),
    .C1(_05433_),
    .C2(_05339_),
    .ZN(_06769_));
 AOI211_X1 _31838_ (.A(_05295_),
    .B(_05342_),
    .C1(_05164_),
    .C2(_05166_),
    .ZN(_06770_));
 NAND4_X1 _31839_ (.A1(_05168_),
    .A2(_05146_),
    .A3(_05438_),
    .A4(_05151_),
    .ZN(_06771_));
 NAND4_X1 _31840_ (.A1(_05438_),
    .A2(_05171_),
    .A3(_05151_),
    .A4(_05172_),
    .ZN(_06772_));
 OAI211_X1 _31841_ (.A(_06771_),
    .B(_06772_),
    .C1(_05342_),
    .C2(_05273_),
    .ZN(_06773_));
 NOR4_X1 _31842_ (.A1(_06769_),
    .A2(_05349_),
    .A3(_06770_),
    .A4(_06773_),
    .ZN(_06774_));
 AOI211_X1 _31843_ (.A(_16682_),
    .B(_05381_),
    .C1(_05140_),
    .C2(_05147_),
    .ZN(_06775_));
 OAI21_X1 _31844_ (.A(_05220_),
    .B1(_05261_),
    .B2(_05177_),
    .ZN(_06777_));
 NAND3_X1 _31845_ (.A1(_05204_),
    .A2(_05220_),
    .A3(_05190_),
    .ZN(_06778_));
 OAI21_X1 _31846_ (.A(_05220_),
    .B1(_05209_),
    .B2(_05332_),
    .ZN(_06779_));
 NAND4_X1 _31847_ (.A1(_06777_),
    .A2(_06778_),
    .A3(_06779_),
    .A4(_06416_),
    .ZN(_06780_));
 OAI211_X1 _31848_ (.A(_05380_),
    .B(_05135_),
    .C1(_05122_),
    .C2(_05165_),
    .ZN(_06781_));
 NAND2_X1 _31849_ (.A1(_05237_),
    .A2(_05380_),
    .ZN(_06782_));
 NAND2_X1 _31850_ (.A1(_06781_),
    .A2(_06782_),
    .ZN(_06783_));
 NOR3_X1 _31851_ (.A1(_06775_),
    .A2(_06780_),
    .A3(_06783_),
    .ZN(_06784_));
 OAI21_X1 _31852_ (.A(_05358_),
    .B1(_05252_),
    .B2(_05301_),
    .ZN(_06785_));
 AND2_X1 _31853_ (.A1(_05329_),
    .A2(_05142_),
    .ZN(_06786_));
 AND2_X1 _31854_ (.A1(_05328_),
    .A2(_05176_),
    .ZN(_06788_));
 AND2_X1 _31855_ (.A1(_05329_),
    .A2(_05316_),
    .ZN(_06789_));
 NOR4_X1 _31856_ (.A1(_06365_),
    .A2(_06786_),
    .A3(_06788_),
    .A4(_06789_),
    .ZN(_06790_));
 OAI21_X1 _31857_ (.A(_05358_),
    .B1(_05312_),
    .B2(_05284_),
    .ZN(_06791_));
 OAI211_X1 _31858_ (.A(_05358_),
    .B(_16682_),
    .C1(_05140_),
    .C2(_05147_),
    .ZN(_06792_));
 AND4_X1 _31859_ (.A1(_06785_),
    .A2(_06790_),
    .A3(_06791_),
    .A4(_06792_),
    .ZN(_06793_));
 AND4_X1 _31860_ (.A1(_06763_),
    .A2(_06774_),
    .A3(_06784_),
    .A4(_06793_),
    .ZN(_06794_));
 AND2_X1 _31861_ (.A1(_05314_),
    .A2(_05321_),
    .ZN(_06795_));
 OAI21_X1 _31862_ (.A(_05297_),
    .B1(_06360_),
    .B2(_05183_),
    .ZN(_06796_));
 OAI21_X1 _31863_ (.A(_05311_),
    .B1(_05462_),
    .B2(_05237_),
    .ZN(_06797_));
 NAND2_X1 _31864_ (.A1(_05297_),
    .A2(_05261_),
    .ZN(_06799_));
 NAND3_X1 _31865_ (.A1(_05219_),
    .A2(_06394_),
    .A3(_06767_),
    .ZN(_06800_));
 AND3_X1 _31866_ (.A1(_05391_),
    .A2(_06799_),
    .A3(_06800_),
    .ZN(_06801_));
 AND4_X1 _31867_ (.A1(_06795_),
    .A2(_06796_),
    .A3(_06797_),
    .A4(_06801_),
    .ZN(_06802_));
 OR2_X1 _31868_ (.A1(_06759_),
    .A2(_06374_),
    .ZN(_06803_));
 NAND4_X1 _31869_ (.A1(_05175_),
    .A2(_05164_),
    .A3(_05172_),
    .A4(_05168_),
    .ZN(_06804_));
 NAND2_X1 _31870_ (.A1(_06803_),
    .A2(_06804_),
    .ZN(_06805_));
 INV_X1 _31871_ (.A(_05398_),
    .ZN(_06806_));
 NAND2_X1 _31872_ (.A1(_05316_),
    .A2(_05187_),
    .ZN(_06807_));
 OAI21_X1 _31873_ (.A(_06384_),
    .B1(_05446_),
    .B2(_05312_),
    .ZN(_06808_));
 NAND4_X1 _31874_ (.A1(_06806_),
    .A2(_05472_),
    .A3(_06807_),
    .A4(_06808_),
    .ZN(_06810_));
 AND2_X1 _31875_ (.A1(_05301_),
    .A2(_05175_),
    .ZN(_06811_));
 AND2_X1 _31876_ (.A1(_05331_),
    .A2(_05175_),
    .ZN(_06812_));
 NOR4_X1 _31877_ (.A1(_06805_),
    .A2(_06810_),
    .A3(_06811_),
    .A4(_06812_),
    .ZN(_06813_));
 OAI21_X1 _31878_ (.A(_05281_),
    .B1(_05219_),
    .B2(_05213_),
    .ZN(_06814_));
 OAI21_X1 _31879_ (.A(_05281_),
    .B1(_05384_),
    .B2(_05332_),
    .ZN(_06815_));
 OAI21_X1 _31880_ (.A(_05441_),
    .B1(_05219_),
    .B2(_05312_),
    .ZN(_06816_));
 OAI21_X1 _31881_ (.A(_05441_),
    .B1(_05384_),
    .B2(_05256_),
    .ZN(_06817_));
 AND4_X1 _31882_ (.A1(_06814_),
    .A2(_06815_),
    .A3(_06816_),
    .A4(_06817_),
    .ZN(_06818_));
 AND2_X1 _31883_ (.A1(_05134_),
    .A2(_05136_),
    .ZN(_06819_));
 OAI21_X1 _31884_ (.A(_05143_),
    .B1(_06819_),
    .B2(_05256_),
    .ZN(_06821_));
 NAND4_X1 _31885_ (.A1(_05151_),
    .A2(_05200_),
    .A3(_05152_),
    .A4(_05140_),
    .ZN(_06822_));
 NAND3_X1 _31886_ (.A1(_05143_),
    .A2(_05201_),
    .A3(_05190_),
    .ZN(_06823_));
 AND3_X1 _31887_ (.A1(_06821_),
    .A2(_06822_),
    .A3(_06823_),
    .ZN(_06824_));
 NAND2_X1 _31888_ (.A1(_05199_),
    .A2(_05127_),
    .ZN(_06825_));
 NAND3_X1 _31889_ (.A1(_05384_),
    .A2(_06767_),
    .A3(_05152_),
    .ZN(_06826_));
 NAND3_X1 _31890_ (.A1(_05462_),
    .A2(_06767_),
    .A3(_05152_),
    .ZN(_06827_));
 AND3_X1 _31891_ (.A1(_06825_),
    .A2(_06826_),
    .A3(_06827_),
    .ZN(_06828_));
 NAND4_X1 _31892_ (.A1(_06767_),
    .A2(_05124_),
    .A3(_05200_),
    .A4(_05152_),
    .ZN(_06829_));
 AND2_X1 _31893_ (.A1(_05425_),
    .A2(_06829_),
    .ZN(_06830_));
 OAI21_X1 _31894_ (.A(_05199_),
    .B1(_05252_),
    .B2(_05301_),
    .ZN(_06832_));
 AND4_X1 _31895_ (.A1(_06824_),
    .A2(_06828_),
    .A3(_06830_),
    .A4(_06832_),
    .ZN(_06833_));
 AND4_X1 _31896_ (.A1(_06802_),
    .A2(_06813_),
    .A3(_06818_),
    .A4(_06833_),
    .ZN(_06834_));
 NAND2_X2 _31897_ (.A1(_06794_),
    .A2(_06834_),
    .ZN(_06835_));
 XOR2_X2 _31898_ (.A(_06757_),
    .B(_06835_),
    .Z(_06836_));
 INV_X1 _31899_ (.A(_06156_),
    .ZN(_06837_));
 NAND2_X1 _31900_ (.A1(_06153_),
    .A2(_06101_),
    .ZN(_06838_));
 NAND3_X1 _31901_ (.A1(_06837_),
    .A2(_06152_),
    .A3(_06838_),
    .ZN(_06839_));
 AND2_X1 _31902_ (.A1(_06033_),
    .A2(_06153_),
    .ZN(_06840_));
 NAND2_X1 _31903_ (.A1(_06153_),
    .A2(_06107_),
    .ZN(_06841_));
 NAND2_X1 _31904_ (.A1(_06157_),
    .A2(_06841_),
    .ZN(_06843_));
 CLKBUF_X2 _31905_ (.A(_06180_),
    .Z(_06844_));
 NAND2_X1 _31906_ (.A1(_06844_),
    .A2(_06107_),
    .ZN(_06845_));
 NAND2_X1 _31907_ (.A1(_06180_),
    .A2(_06099_),
    .ZN(_06846_));
 NAND4_X1 _31908_ (.A1(_06845_),
    .A2(_06187_),
    .A3(_06189_),
    .A4(_06846_),
    .ZN(_06847_));
 NOR4_X1 _31909_ (.A1(_06839_),
    .A2(_06840_),
    .A3(_06843_),
    .A4(_06847_),
    .ZN(_06848_));
 BUF_X2 _31910_ (.A(_06038_),
    .Z(_06849_));
 OAI21_X1 _31911_ (.A(_06849_),
    .B1(_06521_),
    .B2(_06170_),
    .ZN(_06850_));
 INV_X2 _31912_ (.A(_06143_),
    .ZN(_06851_));
 AOI21_X1 _31913_ (.A(_06064_),
    .B1(_06042_),
    .B2(_06851_),
    .ZN(_06852_));
 AND4_X1 _31914_ (.A1(_06009_),
    .A2(_06059_),
    .A3(_06183_),
    .A4(_05993_),
    .ZN(_06854_));
 NOR3_X1 _31915_ (.A1(_06852_),
    .A2(_06070_),
    .A3(_06854_),
    .ZN(_06855_));
 NAND2_X1 _31916_ (.A1(_06849_),
    .A2(_06177_),
    .ZN(_06856_));
 OAI21_X1 _31917_ (.A(_06849_),
    .B1(_06168_),
    .B2(_06128_),
    .ZN(_06857_));
 AND4_X1 _31918_ (.A1(_06850_),
    .A2(_06855_),
    .A3(_06856_),
    .A4(_06857_),
    .ZN(_06858_));
 OAI21_X1 _31919_ (.A(_06137_),
    .B1(_06101_),
    .B2(_06103_),
    .ZN(_06859_));
 BUF_X2 _31920_ (.A(_06163_),
    .Z(_06860_));
 OAI21_X1 _31921_ (.A(_06167_),
    .B1(_06101_),
    .B2(_06860_),
    .ZN(_06861_));
 OAI21_X1 _31922_ (.A(_06167_),
    .B1(_06091_),
    .B2(_06130_),
    .ZN(_06862_));
 OAI21_X1 _31923_ (.A(_06137_),
    .B1(_06091_),
    .B2(_06049_),
    .ZN(_06863_));
 AND4_X1 _31924_ (.A1(_06859_),
    .A2(_06861_),
    .A3(_06862_),
    .A4(_06863_),
    .ZN(_06865_));
 INV_X1 _31925_ (.A(_05997_),
    .ZN(_06866_));
 NOR2_X1 _31926_ (.A1(_06866_),
    .A2(_06509_),
    .ZN(_06867_));
 NOR2_X1 _31927_ (.A1(_06867_),
    .A2(_06488_),
    .ZN(_06868_));
 AND2_X1 _31928_ (.A1(_06027_),
    .A2(_06013_),
    .ZN(_06869_));
 NAND2_X1 _31929_ (.A1(_06023_),
    .A2(_06869_),
    .ZN(_06870_));
 INV_X1 _31930_ (.A(_06023_),
    .ZN(_06871_));
 INV_X1 _31931_ (.A(_06069_),
    .ZN(_06872_));
 OAI21_X1 _31932_ (.A(_06870_),
    .B1(_06871_),
    .B2(_06872_),
    .ZN(_06873_));
 AND3_X1 _31933_ (.A1(_06095_),
    .A2(_06172_),
    .A3(_05993_),
    .ZN(_06874_));
 AND2_X1 _31934_ (.A1(_06023_),
    .A2(_06211_),
    .ZN(_06876_));
 NOR3_X1 _31935_ (.A1(_06873_),
    .A2(_06874_),
    .A3(_06876_),
    .ZN(_06877_));
 OAI21_X1 _31936_ (.A(_05997_),
    .B1(_06200_),
    .B2(_06168_),
    .ZN(_06878_));
 OAI21_X1 _31937_ (.A(_06035_),
    .B1(_06146_),
    .B2(_06860_),
    .ZN(_06879_));
 AND4_X1 _31938_ (.A1(_06868_),
    .A2(_06877_),
    .A3(_06878_),
    .A4(_06879_),
    .ZN(_06880_));
 AND4_X1 _31939_ (.A1(_06848_),
    .A2(_06858_),
    .A3(_06865_),
    .A4(_06880_),
    .ZN(_06881_));
 OAI21_X1 _31940_ (.A(_06450_),
    .B1(_06458_),
    .B2(_06088_),
    .ZN(_06882_));
 INV_X1 _31941_ (.A(_06522_),
    .ZN(_06883_));
 AOI21_X1 _31942_ (.A(_06120_),
    .B1(_06883_),
    .B2(_06509_),
    .ZN(_06884_));
 INV_X1 _31943_ (.A(_06130_),
    .ZN(_06885_));
 AOI21_X1 _31944_ (.A(_06088_),
    .B1(_06514_),
    .B2(_06885_),
    .ZN(_06887_));
 NOR4_X1 _31945_ (.A1(_06882_),
    .A2(_06884_),
    .A3(_06445_),
    .A4(_06887_),
    .ZN(_06888_));
 CLKBUF_X2 _31946_ (.A(_06211_),
    .Z(_06889_));
 NAND2_X1 _31947_ (.A1(_06224_),
    .A2(_06889_),
    .ZN(_06890_));
 AND2_X1 _31948_ (.A1(_06196_),
    .A2(_06000_),
    .ZN(_06891_));
 INV_X1 _31949_ (.A(_06891_),
    .ZN(_06892_));
 NAND2_X1 _31950_ (.A1(_06197_),
    .A2(_06211_),
    .ZN(_06893_));
 NAND3_X1 _31951_ (.A1(_06095_),
    .A2(_06172_),
    .A3(_06213_),
    .ZN(_06894_));
 AND4_X1 _31952_ (.A1(_06892_),
    .A2(_06549_),
    .A3(_06893_),
    .A4(_06894_),
    .ZN(_06895_));
 AND2_X1 _31953_ (.A1(_06221_),
    .A2(_06177_),
    .ZN(_06896_));
 AOI211_X1 _31954_ (.A(_06896_),
    .B(_06222_),
    .C1(_06168_),
    .C2(_06224_),
    .ZN(_06898_));
 OAI21_X1 _31955_ (.A(_06224_),
    .B1(_06099_),
    .B2(_06482_),
    .ZN(_06899_));
 AND4_X1 _31956_ (.A1(_06890_),
    .A2(_06895_),
    .A3(_06898_),
    .A4(_06899_),
    .ZN(_06900_));
 AND2_X1 _31957_ (.A1(_06097_),
    .A2(_06048_),
    .ZN(_06901_));
 INV_X1 _31958_ (.A(_06901_),
    .ZN(_06902_));
 OAI211_X1 _31959_ (.A(_06902_),
    .B(_06472_),
    .C1(_06883_),
    .C2(_06464_),
    .ZN(_06903_));
 AND3_X1 _31960_ (.A1(_06090_),
    .A2(_16760_),
    .A3(_06011_),
    .ZN(_06904_));
 AND2_X1 _31961_ (.A1(_06097_),
    .A2(_06075_),
    .ZN(_06905_));
 OR2_X1 _31962_ (.A1(_06904_),
    .A2(_06905_),
    .ZN(_06906_));
 OAI21_X1 _31963_ (.A(_06111_),
    .B1(_06107_),
    .B2(_06114_),
    .ZN(_06907_));
 NAND2_X1 _31964_ (.A1(_06091_),
    .A2(_06111_),
    .ZN(_06909_));
 NAND2_X1 _31965_ (.A1(_06907_),
    .A2(_06909_),
    .ZN(_06910_));
 NAND3_X1 _31966_ (.A1(_06111_),
    .A2(_06007_),
    .A3(_06198_),
    .ZN(_06911_));
 NAND2_X1 _31967_ (.A1(_06080_),
    .A2(_06110_),
    .ZN(_06912_));
 NAND3_X1 _31968_ (.A1(_06110_),
    .A2(_06008_),
    .A3(_06007_),
    .ZN(_06913_));
 NAND2_X1 _31969_ (.A1(_06110_),
    .A2(_06000_),
    .ZN(_06914_));
 NAND4_X1 _31970_ (.A1(_06911_),
    .A2(_06912_),
    .A3(_06913_),
    .A4(_06914_),
    .ZN(_06915_));
 NOR4_X1 _31971_ (.A1(_06903_),
    .A2(_06906_),
    .A3(_06910_),
    .A4(_06915_),
    .ZN(_06916_));
 OAI211_X1 _31972_ (.A(_06202_),
    .B(_06005_),
    .C1(_06044_),
    .C2(_06045_),
    .ZN(_06917_));
 OAI211_X1 _31973_ (.A(_06202_),
    .B(_06014_),
    .C1(_06044_),
    .C2(_06045_),
    .ZN(_06918_));
 OAI21_X1 _31974_ (.A(_06202_),
    .B1(_06086_),
    .B2(_06052_),
    .ZN(_06920_));
 AND4_X1 _31975_ (.A1(_06203_),
    .A2(_06917_),
    .A3(_06918_),
    .A4(_06920_),
    .ZN(_06921_));
 OAI211_X1 _31976_ (.A(_06210_),
    .B(_06007_),
    .C1(_06032_),
    .C2(_06150_),
    .ZN(_06922_));
 NOR2_X1 _31977_ (.A1(_05989_),
    .A2(_06150_),
    .ZN(_06923_));
 OAI21_X1 _31978_ (.A(_06210_),
    .B1(_06923_),
    .B2(_06091_),
    .ZN(_06924_));
 AND4_X1 _31979_ (.A1(_06530_),
    .A2(_06921_),
    .A3(_06922_),
    .A4(_06924_),
    .ZN(_06925_));
 AND4_X1 _31980_ (.A1(_06888_),
    .A2(_06900_),
    .A3(_06916_),
    .A4(_06925_),
    .ZN(_06926_));
 AND2_X2 _31981_ (.A1(_06881_),
    .A2(_06926_),
    .ZN(_06927_));
 XNOR2_X1 _31982_ (.A(_06927_),
    .B(_00991_),
    .ZN(_06928_));
 XNOR2_X1 _31983_ (.A(_06836_),
    .B(_06928_),
    .ZN(_06929_));
 OAI21_X1 _31984_ (.A(_05957_),
    .B1(_05846_),
    .B2(_05783_),
    .ZN(_06931_));
 NAND2_X1 _31985_ (.A1(_05744_),
    .A2(_05957_),
    .ZN(_06932_));
 NAND4_X1 _31986_ (.A1(_05948_),
    .A2(_05887_),
    .A3(_05759_),
    .A4(_05748_),
    .ZN(_06933_));
 NAND3_X1 _31987_ (.A1(_06931_),
    .A2(_06932_),
    .A3(_06933_),
    .ZN(_06934_));
 AND3_X1 _31988_ (.A1(_05854_),
    .A2(_05947_),
    .A3(_05825_),
    .ZN(_06935_));
 AND2_X1 _31989_ (.A1(_05972_),
    .A2(_05862_),
    .ZN(_06936_));
 AND2_X1 _31990_ (.A1(_05972_),
    .A2(_06660_),
    .ZN(_06937_));
 AND2_X1 _31991_ (.A1(_05972_),
    .A2(_05831_),
    .ZN(_06938_));
 OR4_X1 _31992_ (.A1(_06935_),
    .A2(_06936_),
    .A3(_06937_),
    .A4(_06938_),
    .ZN(_06939_));
 AND2_X1 _31993_ (.A1(_05952_),
    .A2(_05778_),
    .ZN(_06940_));
 AND2_X1 _31994_ (.A1(_05952_),
    .A2(_05811_),
    .ZN(_06942_));
 AND2_X1 _31995_ (.A1(_05950_),
    .A2(_05788_),
    .ZN(_06943_));
 AND3_X1 _31996_ (.A1(_05773_),
    .A2(_05756_),
    .A3(_05947_),
    .ZN(_06944_));
 OR4_X1 _31997_ (.A1(_06940_),
    .A2(_06942_),
    .A3(_06943_),
    .A4(_06944_),
    .ZN(_06945_));
 OAI21_X1 _31998_ (.A(_05967_),
    .B1(_06605_),
    .B2(_06595_),
    .ZN(_06946_));
 NAND3_X1 _31999_ (.A1(_06570_),
    .A2(_05948_),
    .A3(_05802_),
    .ZN(_06947_));
 INV_X1 _32000_ (.A(_05856_),
    .ZN(_06948_));
 OAI211_X1 _32001_ (.A(_06946_),
    .B(_06947_),
    .C1(_06948_),
    .C2(_06591_),
    .ZN(_06949_));
 OR4_X1 _32002_ (.A1(_06934_),
    .A2(_06939_),
    .A3(_06945_),
    .A4(_06949_),
    .ZN(_06950_));
 OAI21_X1 _32003_ (.A(_05909_),
    .B1(_05931_),
    .B2(_05837_),
    .ZN(_06951_));
 AND2_X1 _32004_ (.A1(_05816_),
    .A2(_05899_),
    .ZN(_06953_));
 AND2_X1 _32005_ (.A1(_05788_),
    .A2(_05898_),
    .ZN(_06954_));
 NOR4_X1 _32006_ (.A1(_05919_),
    .A2(_06953_),
    .A3(_06954_),
    .A4(_05920_),
    .ZN(_06955_));
 NAND2_X1 _32007_ (.A1(_05856_),
    .A2(_05899_),
    .ZN(_06956_));
 OAI211_X1 _32008_ (.A(_05908_),
    .B(_05739_),
    .C1(_05745_),
    .C2(_05781_),
    .ZN(_06957_));
 AND4_X1 _32009_ (.A1(_06951_),
    .A2(_06955_),
    .A3(_06956_),
    .A4(_06957_),
    .ZN(_06958_));
 NAND3_X1 _32010_ (.A1(_06604_),
    .A2(_05821_),
    .A3(_06582_),
    .ZN(_06959_));
 INV_X1 _32011_ (.A(_05938_),
    .ZN(_06960_));
 INV_X1 _32012_ (.A(_06618_),
    .ZN(_06961_));
 AOI21_X1 _32013_ (.A(_06960_),
    .B1(_06599_),
    .B2(_06961_),
    .ZN(_06962_));
 AND2_X1 _32014_ (.A1(_06559_),
    .A2(_05938_),
    .ZN(_06964_));
 AND2_X1 _32015_ (.A1(_05930_),
    .A2(_05938_),
    .ZN(_06965_));
 NOR4_X1 _32016_ (.A1(_06962_),
    .A2(_05944_),
    .A3(_06964_),
    .A4(_06965_),
    .ZN(_06966_));
 OAI21_X1 _32017_ (.A(_06604_),
    .B1(_05955_),
    .B2(_05817_),
    .ZN(_06967_));
 NAND4_X1 _32018_ (.A1(_06958_),
    .A2(_06959_),
    .A3(_06966_),
    .A4(_06967_),
    .ZN(_06968_));
 INV_X1 _32019_ (.A(_05826_),
    .ZN(_06969_));
 INV_X1 _32020_ (.A(_05969_),
    .ZN(_06970_));
 AOI21_X1 _32021_ (.A(_06969_),
    .B1(_05889_),
    .B2(_06970_),
    .ZN(_06971_));
 AND2_X1 _32022_ (.A1(_05826_),
    .A2(_05862_),
    .ZN(_06972_));
 AND2_X1 _32023_ (.A1(_05826_),
    .A2(_05831_),
    .ZN(_06973_));
 NOR2_X1 _32024_ (.A1(_06972_),
    .A2(_06973_),
    .ZN(_06975_));
 INV_X1 _32025_ (.A(_06975_),
    .ZN(_06976_));
 AND2_X1 _32026_ (.A1(_05739_),
    .A2(_05745_),
    .ZN(_06977_));
 AOI211_X1 _32027_ (.A(_06971_),
    .B(_06976_),
    .C1(_06977_),
    .C2(_05827_),
    .ZN(_06978_));
 OAI21_X1 _32028_ (.A(_05860_),
    .B1(_06605_),
    .B2(_05804_),
    .ZN(_06979_));
 AND2_X1 _32029_ (.A1(_05860_),
    .A2(_05833_),
    .ZN(_06980_));
 INV_X1 _32030_ (.A(_06980_),
    .ZN(_06981_));
 INV_X1 _32031_ (.A(_06607_),
    .ZN(_06982_));
 NAND2_X1 _32032_ (.A1(_06982_),
    .A2(_05860_),
    .ZN(_06983_));
 AND3_X1 _32033_ (.A1(_06979_),
    .A2(_06981_),
    .A3(_06983_),
    .ZN(_06984_));
 NAND2_X1 _32034_ (.A1(_05842_),
    .A2(_05817_),
    .ZN(_06986_));
 INV_X1 _32035_ (.A(_05788_),
    .ZN(_06987_));
 OAI21_X1 _32036_ (.A(_06986_),
    .B1(_06643_),
    .B2(_06987_),
    .ZN(_06988_));
 AOI21_X1 _32037_ (.A(_06643_),
    .B1(_05961_),
    .B2(_05769_),
    .ZN(_06989_));
 AOI211_X1 _32038_ (.A(_06988_),
    .B(_06989_),
    .C1(_05955_),
    .C2(_05843_),
    .ZN(_06990_));
 AND4_X1 _32039_ (.A1(_05872_),
    .A2(_05844_),
    .A3(_05849_),
    .A4(_05802_),
    .ZN(_06991_));
 AND4_X1 _32040_ (.A1(_05763_),
    .A2(_05739_),
    .A3(_05849_),
    .A4(_05802_),
    .ZN(_06992_));
 NOR4_X1 _32041_ (.A1(_05824_),
    .A2(_06991_),
    .A3(_05805_),
    .A4(_06992_),
    .ZN(_06993_));
 NAND4_X1 _32042_ (.A1(_06978_),
    .A2(_06984_),
    .A3(_06990_),
    .A4(_06993_),
    .ZN(_06994_));
 NOR2_X1 _32043_ (.A1(_05871_),
    .A2(_06607_),
    .ZN(_06995_));
 INV_X1 _32044_ (.A(_05773_),
    .ZN(_06997_));
 AOI21_X1 _32045_ (.A(_05871_),
    .B1(_06997_),
    .B2(_05960_),
    .ZN(_06998_));
 AOI211_X1 _32046_ (.A(_06995_),
    .B(_06998_),
    .C1(_06561_),
    .C2(_05937_),
    .ZN(_06999_));
 NAND2_X1 _32047_ (.A1(_05757_),
    .A2(_05969_),
    .ZN(_07000_));
 NAND2_X1 _32048_ (.A1(_05793_),
    .A2(_07000_),
    .ZN(_07001_));
 AOI211_X1 _32049_ (.A(_05761_),
    .B(_07001_),
    .C1(_06977_),
    .C2(_05771_),
    .ZN(_07002_));
 AND3_X1 _32050_ (.A1(_05750_),
    .A2(_05872_),
    .A3(_05739_),
    .ZN(_07003_));
 AND2_X1 _32051_ (.A1(_05750_),
    .A2(_05831_),
    .ZN(_07004_));
 AND2_X1 _32052_ (.A1(_05750_),
    .A2(_05778_),
    .ZN(_07005_));
 NOR4_X1 _32053_ (.A1(_06625_),
    .A2(_07003_),
    .A3(_07004_),
    .A4(_07005_),
    .ZN(_07006_));
 OAI21_X1 _32054_ (.A(_05883_),
    .B1(_06575_),
    .B2(_06618_),
    .ZN(_07008_));
 OAI211_X1 _32055_ (.A(_05883_),
    .B(_05833_),
    .C1(_05746_),
    .C2(_05763_),
    .ZN(_07009_));
 NAND2_X1 _32056_ (.A1(_05930_),
    .A2(_05882_),
    .ZN(_07010_));
 OAI211_X1 _32057_ (.A(_05882_),
    .B(_05778_),
    .C1(_05745_),
    .C2(_05781_),
    .ZN(_07011_));
 AND4_X1 _32058_ (.A1(_07008_),
    .A2(_07009_),
    .A3(_07010_),
    .A4(_07011_),
    .ZN(_07012_));
 NAND4_X1 _32059_ (.A1(_06999_),
    .A2(_07002_),
    .A3(_07006_),
    .A4(_07012_),
    .ZN(_07013_));
 NOR4_X1 _32060_ (.A1(_06950_),
    .A2(_06968_),
    .A3(_06994_),
    .A4(_07013_),
    .ZN(_07014_));
 AND2_X1 _32061_ (.A1(_06580_),
    .A2(_06581_),
    .ZN(_07015_));
 INV_X1 _32062_ (.A(_07015_),
    .ZN(_07016_));
 NAND2_X2 _32063_ (.A1(_07014_),
    .A2(_07016_),
    .ZN(_07017_));
 XNOR2_X1 _32064_ (.A(_07017_),
    .B(_06437_),
    .ZN(_07019_));
 XNOR2_X1 _32065_ (.A(_06929_),
    .B(_07019_),
    .ZN(_07020_));
 MUX2_X1 _32066_ (.A(_06674_),
    .B(_07020_),
    .S(_05069_),
    .Z(_00702_));
 MUX2_X1 _32067_ (.A(_16953_),
    .B(_16825_),
    .S(_06673_),
    .Z(_00750_));
 MUX2_X1 _32068_ (.A(_16954_),
    .B(_16826_),
    .S(_06673_),
    .Z(_00751_));
 MUX2_X1 _32069_ (.A(_16955_),
    .B(_16827_),
    .S(_06673_),
    .Z(_00752_));
 MUX2_X1 _32070_ (.A(_16956_),
    .B(_16828_),
    .S(_06673_),
    .Z(_00753_));
 MUX2_X1 _32071_ (.A(_16958_),
    .B(_16830_),
    .S(_06673_),
    .Z(_00755_));
 MUX2_X1 _32072_ (.A(_16959_),
    .B(_16831_),
    .S(_03836_),
    .Z(_00756_));
 MUX2_X1 _32073_ (.A(_16960_),
    .B(_16832_),
    .S(_03836_),
    .Z(_00757_));
 MUX2_X1 _32074_ (.A(_16961_),
    .B(_16833_),
    .S(_03836_),
    .Z(_00758_));
 MUX2_X1 _32075_ (.A(_16962_),
    .B(_16834_),
    .S(_03836_),
    .Z(_00759_));
 MUX2_X1 _32076_ (.A(_16963_),
    .B(_16835_),
    .S(_03836_),
    .Z(_00760_));
 XOR2_X1 _32077_ (.A(_17124_),
    .B(_17061_),
    .Z(_07022_));
 XOR2_X2 _32078_ (.A(_05484_),
    .B(_06835_),
    .Z(_07023_));
 NOR2_X1 _32079_ (.A1(_06117_),
    .A2(_06098_),
    .ZN(_07024_));
 CLKBUF_X2 _32080_ (.A(_06063_),
    .Z(_07025_));
 NOR2_X1 _32081_ (.A1(_06205_),
    .A2(_06198_),
    .ZN(_07026_));
 AOI221_X4 _32082_ (.A(_07024_),
    .B1(_06143_),
    .B2(_06110_),
    .C1(_07025_),
    .C2(_07026_),
    .ZN(_07027_));
 AND2_X1 _32083_ (.A1(_06167_),
    .A2(_06099_),
    .ZN(_07028_));
 INV_X1 _32084_ (.A(_07028_),
    .ZN(_07030_));
 AND2_X1 _32085_ (.A1(_06166_),
    .A2(_06085_),
    .ZN(_07031_));
 INV_X1 _32086_ (.A(_07031_),
    .ZN(_07032_));
 NAND4_X1 _32087_ (.A1(_06172_),
    .A2(_06158_),
    .A3(_06044_),
    .A4(_06058_),
    .ZN(_07033_));
 AND3_X1 _32088_ (.A1(_07032_),
    .A2(_06173_),
    .A3(_07033_),
    .ZN(_07034_));
 AND2_X1 _32089_ (.A1(_06522_),
    .A2(_06197_),
    .ZN(_07035_));
 INV_X1 _32090_ (.A(_07035_),
    .ZN(_07036_));
 NAND3_X1 _32091_ (.A1(_06188_),
    .A2(_06172_),
    .A3(_06213_),
    .ZN(_07037_));
 AND4_X1 _32092_ (.A1(_07030_),
    .A2(_07034_),
    .A3(_07036_),
    .A4(_07037_),
    .ZN(_07038_));
 AND2_X1 _32093_ (.A1(_06035_),
    .A2(_06128_),
    .ZN(_07039_));
 AND2_X1 _32094_ (.A1(_06166_),
    .A2(_06188_),
    .ZN(_07041_));
 AOI211_X1 _32095_ (.A(_07039_),
    .B(_07041_),
    .C1(_06482_),
    .C2(_06167_),
    .ZN(_07042_));
 OAI21_X1 _32096_ (.A(_06137_),
    .B1(_06869_),
    .B2(_06124_),
    .ZN(_07043_));
 AND2_X1 _32097_ (.A1(_06210_),
    .A2(_06151_),
    .ZN(_07044_));
 NOR2_X1 _32098_ (.A1(_06217_),
    .A2(_07044_),
    .ZN(_07045_));
 OAI21_X1 _32099_ (.A(_06097_),
    .B1(_06080_),
    .B2(_06151_),
    .ZN(_07046_));
 NAND2_X1 _32100_ (.A1(_06038_),
    .A2(_06188_),
    .ZN(_07047_));
 AND4_X1 _32101_ (.A1(_07043_),
    .A2(_07045_),
    .A3(_07046_),
    .A4(_07047_),
    .ZN(_07048_));
 AND4_X1 _32102_ (.A1(_07027_),
    .A2(_07038_),
    .A3(_07042_),
    .A4(_07048_),
    .ZN(_07049_));
 AOI21_X1 _32103_ (.A(_06513_),
    .B1(_06019_),
    .B2(_06137_),
    .ZN(_07050_));
 AND2_X1 _32104_ (.A1(_06091_),
    .A2(_06209_),
    .ZN(_07052_));
 AND2_X1 _32105_ (.A1(_06080_),
    .A2(_06111_),
    .ZN(_07053_));
 AND3_X1 _32106_ (.A1(_06211_),
    .A2(_05997_),
    .A3(_06065_),
    .ZN(_07054_));
 NOR4_X1 _32107_ (.A1(_06905_),
    .A2(_07052_),
    .A3(_07053_),
    .A4(_07054_),
    .ZN(_07055_));
 AND2_X1 _32108_ (.A1(_06080_),
    .A2(_06221_),
    .ZN(_07056_));
 OR2_X1 _32109_ (.A1(_07056_),
    .A2(_06081_),
    .ZN(_07057_));
 AND3_X1 _32110_ (.A1(_06122_),
    .A2(_06065_),
    .A3(_06889_),
    .ZN(_07058_));
 AND2_X1 _32111_ (.A1(_06210_),
    .A2(_06170_),
    .ZN(_07059_));
 NOR4_X1 _32112_ (.A1(_07057_),
    .A2(_07058_),
    .A3(_07059_),
    .A4(_06461_),
    .ZN(_07060_));
 AOI21_X1 _32113_ (.A(_06088_),
    .B1(_06506_),
    .B2(_06455_),
    .ZN(_07061_));
 AND2_X1 _32114_ (.A1(_06095_),
    .A2(_06122_),
    .ZN(_07063_));
 AND2_X1 _32115_ (.A1(_06869_),
    .A2(_06082_),
    .ZN(_07064_));
 AND3_X1 _32116_ (.A1(_06052_),
    .A2(_06172_),
    .A3(_05993_),
    .ZN(_07065_));
 NOR4_X1 _32117_ (.A1(_07061_),
    .A2(_07063_),
    .A3(_07064_),
    .A4(_07065_),
    .ZN(_07066_));
 AND4_X1 _32118_ (.A1(_07050_),
    .A2(_07055_),
    .A3(_07060_),
    .A4(_07066_),
    .ZN(_07067_));
 OAI21_X1 _32119_ (.A(_06122_),
    .B1(_06076_),
    .B2(_06049_),
    .ZN(_07068_));
 NOR2_X1 _32120_ (.A1(_06096_),
    .A2(_06901_),
    .ZN(_07069_));
 AND2_X1 _32121_ (.A1(_06013_),
    .A2(_06045_),
    .ZN(_07070_));
 OAI21_X1 _32122_ (.A(_06844_),
    .B1(_06041_),
    .B2(_07070_),
    .ZN(_07071_));
 AND2_X1 _32123_ (.A1(_06023_),
    .A2(_06124_),
    .ZN(_07072_));
 INV_X1 _32124_ (.A(_07072_),
    .ZN(_07074_));
 AND4_X1 _32125_ (.A1(_07068_),
    .A2(_07069_),
    .A3(_07071_),
    .A4(_07074_),
    .ZN(_07075_));
 NAND4_X1 _32126_ (.A1(_06213_),
    .A2(_06009_),
    .A3(_06183_),
    .A4(_06043_),
    .ZN(_07076_));
 AOI21_X1 _32127_ (.A(_06866_),
    .B1(_06042_),
    .B2(_06467_),
    .ZN(_07077_));
 AOI211_X1 _32128_ (.A(_06896_),
    .B(_07077_),
    .C1(_06059_),
    .C2(_06197_),
    .ZN(_07078_));
 AND4_X1 _32129_ (.A1(_06008_),
    .A2(_06213_),
    .A3(_06059_),
    .A4(_06183_),
    .ZN(_07079_));
 AND2_X1 _32130_ (.A1(_06107_),
    .A2(_06202_),
    .ZN(_07080_));
 BUF_X2 _32131_ (.A(_06202_),
    .Z(_07081_));
 AOI211_X1 _32132_ (.A(_07079_),
    .B(_07080_),
    .C1(_06033_),
    .C2(_07081_),
    .ZN(_07082_));
 OAI211_X1 _32133_ (.A(_07081_),
    .B(_06007_),
    .C1(_06008_),
    .C2(_06065_),
    .ZN(_07083_));
 AND4_X1 _32134_ (.A1(_07076_),
    .A2(_07078_),
    .A3(_07082_),
    .A4(_07083_),
    .ZN(_07085_));
 NAND4_X1 _32135_ (.A1(_07049_),
    .A2(_07067_),
    .A3(_07075_),
    .A4(_07085_),
    .ZN(_07086_));
 NAND2_X1 _32136_ (.A1(_06923_),
    .A2(_06224_),
    .ZN(_07087_));
 AND2_X1 _32137_ (.A1(_06166_),
    .A2(_06163_),
    .ZN(_07088_));
 AOI221_X4 _32138_ (.A(_07088_),
    .B1(_06038_),
    .B2(_06076_),
    .C1(_06035_),
    .C2(_06033_),
    .ZN(_07089_));
 AND2_X1 _32139_ (.A1(_06058_),
    .A2(_06045_),
    .ZN(_07090_));
 AOI221_X4 _32140_ (.A(_06489_),
    .B1(_06860_),
    .B2(_06180_),
    .C1(_06137_),
    .C2(_07090_),
    .ZN(_07091_));
 AOI221_X4 _32141_ (.A(_06129_),
    .B1(_06000_),
    .B2(_06082_),
    .C1(_06889_),
    .C2(_06111_),
    .ZN(_07092_));
 AND4_X1 _32142_ (.A1(_07087_),
    .A2(_07089_),
    .A3(_07091_),
    .A4(_07092_),
    .ZN(_07093_));
 AOI22_X1 _32143_ (.A1(_06114_),
    .A2(_06153_),
    .B1(_06482_),
    .B2(_06224_),
    .ZN(_07094_));
 OAI221_X1 _32144_ (.A(_07094_),
    .B1(_06098_),
    .B2(_06120_),
    .C1(_06514_),
    .C2(_06088_),
    .ZN(_07096_));
 NAND2_X1 _32145_ (.A1(_06153_),
    .A2(_06049_),
    .ZN(_07097_));
 NAND2_X1 _32146_ (.A1(_06892_),
    .A2(_07097_),
    .ZN(_07098_));
 NOR4_X1 _32147_ (.A1(_07096_),
    .A2(_07098_),
    .A3(_06453_),
    .A4(_06536_),
    .ZN(_07099_));
 AND3_X1 _32148_ (.A1(_06889_),
    .A2(_07025_),
    .A3(_06065_),
    .ZN(_07100_));
 AND2_X1 _32149_ (.A1(_06038_),
    .A2(_06889_),
    .ZN(_07101_));
 AOI221_X4 _32150_ (.A(_07100_),
    .B1(_06103_),
    .B2(_06122_),
    .C1(_06009_),
    .C2(_07101_),
    .ZN(_07102_));
 AND2_X1 _32151_ (.A1(_06086_),
    .A2(_05996_),
    .ZN(_07103_));
 AOI221_X4 _32152_ (.A(_07103_),
    .B1(_06107_),
    .B2(_06180_),
    .C1(_06086_),
    .C2(_06082_),
    .ZN(_07104_));
 AOI22_X1 _32153_ (.A1(_06146_),
    .A2(_06122_),
    .B1(_06860_),
    .B2(_06111_),
    .ZN(_07105_));
 AND4_X1 _32154_ (.A1(_06841_),
    .A2(_07104_),
    .A3(_06838_),
    .A4(_07105_),
    .ZN(_07107_));
 NAND4_X1 _32155_ (.A1(_07093_),
    .A2(_07099_),
    .A3(_07102_),
    .A4(_07107_),
    .ZN(_07108_));
 NOR2_X2 _32156_ (.A1(_07086_),
    .A2(_07108_),
    .ZN(_07109_));
 XNOR2_X1 _32157_ (.A(_07109_),
    .B(_14440_),
    .ZN(_07110_));
 XNOR2_X1 _32158_ (.A(_07023_),
    .B(_07110_),
    .ZN(_07111_));
 AND2_X1 _32159_ (.A1(_05974_),
    .A2(_05817_),
    .ZN(_07112_));
 INV_X1 _32160_ (.A(_05974_),
    .ZN(_07113_));
 AOI211_X1 _32161_ (.A(_05740_),
    .B(_07113_),
    .C1(_05780_),
    .C2(_05781_),
    .ZN(_07114_));
 AOI211_X1 _32162_ (.A(_07112_),
    .B(_07114_),
    .C1(_05974_),
    .C2(_06605_),
    .ZN(_07115_));
 OAI21_X1 _32163_ (.A(_05979_),
    .B1(_05857_),
    .B2(_05811_),
    .ZN(_07116_));
 AND4_X1 _32164_ (.A1(_05948_),
    .A2(_05977_),
    .A3(_05887_),
    .A4(_05802_),
    .ZN(_07118_));
 AOI21_X1 _32165_ (.A(_06591_),
    .B1(_05954_),
    .B2(_06970_),
    .ZN(_07119_));
 AOI211_X1 _32166_ (.A(_07118_),
    .B(_07119_),
    .C1(_05979_),
    .C2(_05789_),
    .ZN(_07120_));
 NAND4_X1 _32167_ (.A1(_07115_),
    .A2(_06594_),
    .A3(_07116_),
    .A4(_07120_),
    .ZN(_07121_));
 AND2_X1 _32168_ (.A1(_05899_),
    .A2(_05867_),
    .ZN(_07122_));
 OR2_X1 _32169_ (.A1(_05919_),
    .A2(_07122_),
    .ZN(_07123_));
 AND2_X1 _32170_ (.A1(_05811_),
    .A2(_05909_),
    .ZN(_07124_));
 INV_X1 _32171_ (.A(_07124_),
    .ZN(_07125_));
 OAI21_X1 _32172_ (.A(_05912_),
    .B1(_05866_),
    .B2(_05867_),
    .ZN(_07126_));
 OAI211_X1 _32173_ (.A(_07125_),
    .B(_07126_),
    .C1(_06599_),
    .C2(_05922_),
    .ZN(_07127_));
 AND3_X1 _32174_ (.A1(_05900_),
    .A2(_05872_),
    .A3(_05844_),
    .ZN(_07129_));
 OR4_X1 _32175_ (.A1(_07123_),
    .A2(_07127_),
    .A3(_07129_),
    .A4(_05903_),
    .ZN(_07130_));
 AND2_X1 _32176_ (.A1(_05958_),
    .A2(_05892_),
    .ZN(_07131_));
 AND2_X1 _32177_ (.A1(_05952_),
    .A2(_05831_),
    .ZN(_07132_));
 INV_X1 _32178_ (.A(_07132_),
    .ZN(_07133_));
 INV_X1 _32179_ (.A(_06943_),
    .ZN(_07134_));
 NAND2_X1 _32180_ (.A1(_05952_),
    .A2(_05794_),
    .ZN(_07135_));
 NAND3_X1 _32181_ (.A1(_05931_),
    .A2(_05848_),
    .A3(_05948_),
    .ZN(_07136_));
 NAND4_X1 _32182_ (.A1(_07133_),
    .A2(_07134_),
    .A3(_07135_),
    .A4(_07136_),
    .ZN(_07137_));
 AOI211_X1 _32183_ (.A(_05785_),
    .B(_06640_),
    .C1(_06572_),
    .C2(_16801_),
    .ZN(_07138_));
 NAND2_X1 _32184_ (.A1(_06662_),
    .A2(_05851_),
    .ZN(_07140_));
 NOR2_X1 _32185_ (.A1(_06640_),
    .A2(_07140_),
    .ZN(_07141_));
 OR4_X1 _32186_ (.A1(_07131_),
    .A2(_07137_),
    .A3(_07138_),
    .A4(_07141_),
    .ZN(_07142_));
 OAI21_X1 _32187_ (.A(_06604_),
    .B1(_05834_),
    .B2(_05817_),
    .ZN(_07143_));
 OAI21_X1 _32188_ (.A(_05925_),
    .B1(_05864_),
    .B2(_05831_),
    .ZN(_07144_));
 OAI211_X1 _32189_ (.A(_05756_),
    .B(_05906_),
    .C1(_06559_),
    .C2(_06609_),
    .ZN(_07145_));
 NAND3_X1 _32190_ (.A1(_05876_),
    .A2(_05756_),
    .A3(_05906_),
    .ZN(_07146_));
 NAND4_X1 _32191_ (.A1(_07143_),
    .A2(_07144_),
    .A3(_07145_),
    .A4(_07146_),
    .ZN(_07147_));
 OAI21_X1 _32192_ (.A(_05939_),
    .B1(_06595_),
    .B2(_05878_),
    .ZN(_07148_));
 NAND2_X1 _32193_ (.A1(_05817_),
    .A2(_05939_),
    .ZN(_07149_));
 NAND2_X1 _32194_ (.A1(_07148_),
    .A2(_07149_),
    .ZN(_07151_));
 AND2_X1 _32195_ (.A1(_05938_),
    .A2(_05831_),
    .ZN(_07152_));
 OR4_X1 _32196_ (.A1(_05936_),
    .A2(_07147_),
    .A3(_07151_),
    .A4(_07152_),
    .ZN(_07153_));
 NOR4_X1 _32197_ (.A1(_07121_),
    .A2(_07130_),
    .A3(_07142_),
    .A4(_07153_),
    .ZN(_07154_));
 NAND2_X1 _32198_ (.A1(_05747_),
    .A2(_05833_),
    .ZN(_07155_));
 NOR2_X1 _32199_ (.A1(_07155_),
    .A2(_05887_),
    .ZN(_07156_));
 OAI21_X1 _32200_ (.A(_05828_),
    .B1(_07156_),
    .B2(_06605_),
    .ZN(_07157_));
 INV_X1 _32201_ (.A(_06972_),
    .ZN(_07158_));
 AND2_X1 _32202_ (.A1(_05855_),
    .A2(_05827_),
    .ZN(_07159_));
 INV_X1 _32203_ (.A(_07159_),
    .ZN(_07160_));
 NAND4_X1 _32204_ (.A1(_07157_),
    .A2(_05836_),
    .A3(_07158_),
    .A4(_07160_),
    .ZN(_07162_));
 BUF_X2 _32205_ (.A(_05959_),
    .Z(_07163_));
 AND2_X1 _32206_ (.A1(_05809_),
    .A2(_07163_),
    .ZN(_07164_));
 INV_X1 _32207_ (.A(_05878_),
    .ZN(_07165_));
 AOI21_X1 _32208_ (.A(_05813_),
    .B1(_07165_),
    .B2(_06987_),
    .ZN(_07166_));
 NOR4_X1 _32209_ (.A1(_07162_),
    .A2(_06619_),
    .A3(_07164_),
    .A4(_07166_),
    .ZN(_07167_));
 NOR2_X1 _32210_ (.A1(_05871_),
    .A2(_07140_),
    .ZN(_07168_));
 AOI211_X1 _32211_ (.A(_05877_),
    .B(_07168_),
    .C1(_05811_),
    .C2(_06561_),
    .ZN(_07169_));
 AND4_X1 _32212_ (.A1(_05779_),
    .A2(_05825_),
    .A3(_05767_),
    .A4(_05749_),
    .ZN(_07170_));
 AND4_X1 _32213_ (.A1(_05833_),
    .A2(_05887_),
    .A3(_05825_),
    .A4(_05749_),
    .ZN(_07171_));
 AOI211_X1 _32214_ (.A(_07170_),
    .B(_07171_),
    .C1(_06561_),
    .C2(_05789_),
    .ZN(_07173_));
 OAI21_X1 _32215_ (.A(_05886_),
    .B1(_06608_),
    .B2(_05829_),
    .ZN(_07174_));
 OAI21_X1 _32216_ (.A(_05886_),
    .B1(_06568_),
    .B2(_05867_),
    .ZN(_07175_));
 AND4_X1 _32217_ (.A1(_07169_),
    .A2(_07173_),
    .A3(_07174_),
    .A4(_07175_),
    .ZN(_07176_));
 OAI21_X1 _32218_ (.A(_05861_),
    .B1(_05855_),
    .B2(_05773_),
    .ZN(_07177_));
 OAI21_X1 _32219_ (.A(_05843_),
    .B1(_05855_),
    .B2(_07163_),
    .ZN(_07178_));
 OAI21_X1 _32220_ (.A(_05843_),
    .B1(_05817_),
    .B2(_05867_),
    .ZN(_07179_));
 OAI21_X1 _32221_ (.A(_05861_),
    .B1(_05817_),
    .B2(_06609_),
    .ZN(_07180_));
 AND4_X1 _32222_ (.A1(_07177_),
    .A2(_07178_),
    .A3(_07179_),
    .A4(_07180_),
    .ZN(_07181_));
 NAND2_X1 _32223_ (.A1(_05876_),
    .A2(_05751_),
    .ZN(_07182_));
 OAI21_X1 _32224_ (.A(_05774_),
    .B1(_05857_),
    .B2(_05959_),
    .ZN(_07184_));
 NAND2_X1 _32225_ (.A1(_05774_),
    .A2(_05931_),
    .ZN(_07185_));
 AND4_X1 _32226_ (.A1(_05790_),
    .A2(_07184_),
    .A3(_05795_),
    .A4(_07185_),
    .ZN(_07186_));
 AND2_X1 _32227_ (.A1(_07005_),
    .A2(_06662_),
    .ZN(_07187_));
 AND3_X1 _32228_ (.A1(_05750_),
    .A2(_05833_),
    .A3(_05887_),
    .ZN(_07188_));
 NOR2_X1 _32229_ (.A1(_07187_),
    .A2(_07188_),
    .ZN(_07189_));
 NAND3_X1 _32230_ (.A1(_06575_),
    .A2(_05872_),
    .A3(_05751_),
    .ZN(_07190_));
 AND4_X1 _32231_ (.A1(_07182_),
    .A2(_07186_),
    .A3(_07189_),
    .A4(_07190_),
    .ZN(_07191_));
 AND4_X1 _32232_ (.A1(_07167_),
    .A2(_07176_),
    .A3(_07181_),
    .A4(_07191_),
    .ZN(_07192_));
 NAND2_X2 _32233_ (.A1(_07154_),
    .A2(_07192_),
    .ZN(_07193_));
 XNOR2_X1 _32234_ (.A(_07193_),
    .B(_05983_),
    .ZN(_07195_));
 OAI21_X1 _32235_ (.A(_05380_),
    .B1(_05312_),
    .B2(_05284_),
    .ZN(_07196_));
 OAI21_X1 _32236_ (.A(_07196_),
    .B1(_05337_),
    .B2(_05381_),
    .ZN(_07197_));
 OAI21_X1 _32237_ (.A(_05220_),
    .B1(_05407_),
    .B2(_05261_),
    .ZN(_07198_));
 INV_X1 _32238_ (.A(_05207_),
    .ZN(_07199_));
 OAI211_X1 _32239_ (.A(_07198_),
    .B(_05386_),
    .C1(_07199_),
    .C2(_05239_),
    .ZN(_07200_));
 OR2_X1 _32240_ (.A1(_05466_),
    .A2(_05226_),
    .ZN(_07201_));
 OAI21_X1 _32241_ (.A(_06426_),
    .B1(_05273_),
    .B2(_05381_),
    .ZN(_07202_));
 OR4_X1 _32242_ (.A1(_07197_),
    .A2(_07200_),
    .A3(_07201_),
    .A4(_07202_),
    .ZN(_07203_));
 OAI21_X1 _32243_ (.A(_05358_),
    .B1(_06360_),
    .B2(_06372_),
    .ZN(_07204_));
 NAND4_X1 _32244_ (.A1(_06410_),
    .A2(_05438_),
    .A3(_05138_),
    .A4(_05227_),
    .ZN(_07206_));
 AND3_X1 _32245_ (.A1(_07204_),
    .A2(_06791_),
    .A3(_07206_),
    .ZN(_07207_));
 AND2_X1 _32246_ (.A1(_05329_),
    .A2(_05320_),
    .ZN(_07208_));
 NOR4_X1 _32247_ (.A1(_05431_),
    .A2(_06368_),
    .A3(_06788_),
    .A4(_07208_),
    .ZN(_07209_));
 NAND4_X1 _32248_ (.A1(_05438_),
    .A2(_05166_),
    .A3(_05151_),
    .A4(_05200_),
    .ZN(_07210_));
 NAND4_X1 _32249_ (.A1(_06410_),
    .A2(_05438_),
    .A3(_05138_),
    .A4(_05151_),
    .ZN(_07211_));
 OAI211_X1 _32250_ (.A(_07210_),
    .B(_07211_),
    .C1(_05433_),
    .C2(_05342_),
    .ZN(_07212_));
 AOI21_X1 _32251_ (.A(_05342_),
    .B1(_07199_),
    .B2(_05378_),
    .ZN(_07213_));
 AND3_X1 _32252_ (.A1(_05180_),
    .A2(_05347_),
    .A3(_05182_),
    .ZN(_07214_));
 NOR3_X1 _32253_ (.A1(_07212_),
    .A2(_07213_),
    .A3(_07214_),
    .ZN(_07215_));
 NAND2_X1 _32254_ (.A1(_06354_),
    .A2(_05389_),
    .ZN(_07217_));
 OAI21_X1 _32255_ (.A(_07217_),
    .B1(_05339_),
    .B2(_05337_),
    .ZN(_07218_));
 AND2_X1 _32256_ (.A1(_06354_),
    .A2(_05127_),
    .ZN(_07219_));
 NOR4_X1 _32257_ (.A1(_07218_),
    .A2(_06764_),
    .A3(_07219_),
    .A4(_06357_),
    .ZN(_07220_));
 NAND4_X1 _32258_ (.A1(_07207_),
    .A2(_07209_),
    .A3(_07215_),
    .A4(_07220_),
    .ZN(_07221_));
 OAI211_X1 _32259_ (.A(_05263_),
    .B(_05168_),
    .C1(_05164_),
    .C2(_05166_),
    .ZN(_07222_));
 OAI211_X1 _32260_ (.A(_05263_),
    .B(_06410_),
    .C1(_05124_),
    .C2(_05138_),
    .ZN(_07223_));
 OAI21_X1 _32261_ (.A(_05263_),
    .B1(_05248_),
    .B2(_05177_),
    .ZN(_07224_));
 NAND4_X1 _32262_ (.A1(_07222_),
    .A2(_07223_),
    .A3(_05272_),
    .A4(_07224_),
    .ZN(_07225_));
 OAI21_X1 _32263_ (.A(_05244_),
    .B1(_05462_),
    .B2(_05316_),
    .ZN(_07226_));
 OAI21_X1 _32264_ (.A(_05244_),
    .B1(_05261_),
    .B2(_05213_),
    .ZN(_07228_));
 OAI21_X1 _32265_ (.A(_05244_),
    .B1(_05446_),
    .B2(_05252_),
    .ZN(_07229_));
 OAI211_X1 _32266_ (.A(_06767_),
    .B(_05267_),
    .C1(_05332_),
    .C2(_05209_),
    .ZN(_07230_));
 NAND4_X1 _32267_ (.A1(_07226_),
    .A2(_07228_),
    .A3(_07229_),
    .A4(_07230_),
    .ZN(_07231_));
 NOR4_X1 _32268_ (.A1(_07203_),
    .A2(_07221_),
    .A3(_07225_),
    .A4(_07231_),
    .ZN(_07232_));
 OAI211_X1 _32269_ (.A(_06394_),
    .B(_06767_),
    .C1(_05237_),
    .C2(_05332_),
    .ZN(_07233_));
 NAND2_X1 _32270_ (.A1(_05297_),
    .A2(_05306_),
    .ZN(_07234_));
 NAND4_X1 _32271_ (.A1(_06407_),
    .A2(_07233_),
    .A3(_06800_),
    .A4(_07234_),
    .ZN(_07235_));
 AOI21_X1 _32272_ (.A(_05393_),
    .B1(_05194_),
    .B2(_05246_),
    .ZN(_07236_));
 AND2_X1 _32273_ (.A1(_05135_),
    .A2(_05172_),
    .ZN(_07237_));
 INV_X1 _32274_ (.A(_07237_),
    .ZN(_07239_));
 AOI21_X1 _32275_ (.A(_05393_),
    .B1(_07239_),
    .B2(_05378_),
    .ZN(_07240_));
 NOR3_X1 _32276_ (.A1(_07235_),
    .A2(_07236_),
    .A3(_07240_),
    .ZN(_07241_));
 NAND2_X1 _32277_ (.A1(_06819_),
    .A2(_05187_),
    .ZN(_07242_));
 NAND3_X1 _32278_ (.A1(_05209_),
    .A2(_05215_),
    .A3(_05152_),
    .ZN(_07243_));
 AND3_X1 _32279_ (.A1(_07242_),
    .A2(_06807_),
    .A3(_07243_),
    .ZN(_07244_));
 OAI21_X1 _32280_ (.A(_06384_),
    .B1(_05248_),
    .B2(_05177_),
    .ZN(_07245_));
 OAI211_X1 _32281_ (.A(_07244_),
    .B(_07245_),
    .C1(_05477_),
    .C2(_05195_),
    .ZN(_07246_));
 OAI21_X1 _32282_ (.A(_05199_),
    .B1(_05261_),
    .B2(_05320_),
    .ZN(_07247_));
 OAI21_X1 _32283_ (.A(_05143_),
    .B1(_05265_),
    .B2(_05389_),
    .ZN(_07248_));
 NAND2_X1 _32284_ (.A1(_05209_),
    .A2(_05143_),
    .ZN(_07250_));
 NAND4_X1 _32285_ (.A1(_07247_),
    .A2(_07248_),
    .A3(_07250_),
    .A4(_05375_),
    .ZN(_07251_));
 NAND3_X1 _32286_ (.A1(_05175_),
    .A2(_05173_),
    .A3(_06410_),
    .ZN(_07252_));
 NAND3_X1 _32287_ (.A1(_05175_),
    .A2(_05146_),
    .A3(_06410_),
    .ZN(_07253_));
 OAI211_X1 _32288_ (.A(_07252_),
    .B(_07253_),
    .C1(_05294_),
    .C2(_06374_),
    .ZN(_07254_));
 NAND2_X1 _32289_ (.A1(_05209_),
    .A2(_05163_),
    .ZN(_07255_));
 NAND4_X1 _32290_ (.A1(_05168_),
    .A2(_05124_),
    .A3(_05227_),
    .A4(_05152_),
    .ZN(_07256_));
 OAI211_X1 _32291_ (.A(_07255_),
    .B(_07256_),
    .C1(_06386_),
    .C2(_06374_),
    .ZN(_07257_));
 NOR4_X1 _32292_ (.A1(_07246_),
    .A2(_07251_),
    .A3(_07254_),
    .A4(_07257_),
    .ZN(_07258_));
 OAI21_X1 _32293_ (.A(_05281_),
    .B1(_05370_),
    .B2(_05414_),
    .ZN(_07259_));
 OAI211_X1 _32294_ (.A(_06394_),
    .B(_05227_),
    .C1(_05248_),
    .C2(_05177_),
    .ZN(_07261_));
 AND3_X1 _32295_ (.A1(_07259_),
    .A2(_06398_),
    .A3(_07261_),
    .ZN(_07262_));
 INV_X1 _32296_ (.A(_05441_),
    .ZN(_07263_));
 OAI21_X1 _32297_ (.A(_06403_),
    .B1(_07263_),
    .B2(_05454_),
    .ZN(_07264_));
 AND2_X1 _32298_ (.A1(_05441_),
    .A2(_05320_),
    .ZN(_07265_));
 AND3_X1 _32299_ (.A1(_05286_),
    .A2(_05215_),
    .A3(_05171_),
    .ZN(_07266_));
 NOR4_X1 _32300_ (.A1(_07264_),
    .A2(_05304_),
    .A3(_07265_),
    .A4(_07266_),
    .ZN(_07267_));
 AND4_X1 _32301_ (.A1(_07241_),
    .A2(_07258_),
    .A3(_07262_),
    .A4(_07267_),
    .ZN(_07268_));
 NAND2_X2 _32302_ (.A1(_07232_),
    .A2(_07268_),
    .ZN(_07269_));
 NOR2_X1 _32303_ (.A1(_06692_),
    .A2(_05652_),
    .ZN(_07270_));
 AOI21_X1 _32304_ (.A(_07270_),
    .B1(_05703_),
    .B2(_05651_),
    .ZN(_07272_));
 NAND4_X1 _32305_ (.A1(_06312_),
    .A2(_06291_),
    .A3(_05572_),
    .A4(_05716_),
    .ZN(_07273_));
 NAND3_X1 _32306_ (.A1(_07272_),
    .A2(_06683_),
    .A3(_07273_),
    .ZN(_07274_));
 AND2_X1 _32307_ (.A1(_06697_),
    .A2(_05642_),
    .ZN(_07275_));
 AOI21_X1 _32308_ (.A(_05649_),
    .B1(_06335_),
    .B2(_06261_),
    .ZN(_07276_));
 NOR4_X1 _32309_ (.A1(_07274_),
    .A2(_07275_),
    .A3(_06299_),
    .A4(_07276_),
    .ZN(_07277_));
 AND4_X1 _32310_ (.A1(_05611_),
    .A2(_06312_),
    .A3(_05715_),
    .A4(_06309_),
    .ZN(_07278_));
 AND4_X1 _32311_ (.A1(_05525_),
    .A2(_06312_),
    .A3(_05572_),
    .A4(_06309_),
    .ZN(_07279_));
 AOI211_X1 _32312_ (.A(_07278_),
    .B(_07279_),
    .C1(_05670_),
    .C2(_05521_),
    .ZN(_07280_));
 AND3_X1 _32313_ (.A1(_05628_),
    .A2(_06309_),
    .A3(_06312_),
    .ZN(_07281_));
 AND4_X1 _32314_ (.A1(_06285_),
    .A2(_05662_),
    .A3(_05657_),
    .A4(_05666_),
    .ZN(_07283_));
 AOI211_X1 _32315_ (.A(_07281_),
    .B(_07283_),
    .C1(_06346_),
    .C2(_05670_),
    .ZN(_07284_));
 AND2_X1 _32316_ (.A1(_05672_),
    .A2(_06267_),
    .ZN(_07285_));
 AOI211_X1 _32317_ (.A(_05675_),
    .B(_07285_),
    .C1(_05543_),
    .C2(_05673_),
    .ZN(_07286_));
 OAI21_X1 _32318_ (.A(_05673_),
    .B1(_06275_),
    .B2(_05570_),
    .ZN(_07287_));
 AND4_X1 _32319_ (.A1(_07280_),
    .A2(_07284_),
    .A3(_07286_),
    .A4(_07287_),
    .ZN(_07288_));
 AND4_X1 _32320_ (.A1(_05714_),
    .A2(_05525_),
    .A3(_05572_),
    .A4(_05716_),
    .ZN(_07289_));
 AND2_X1 _32321_ (.A1(_05619_),
    .A2(_05710_),
    .ZN(_07290_));
 AOI211_X1 _32322_ (.A(_07289_),
    .B(_07290_),
    .C1(_06711_),
    .C2(_05616_),
    .ZN(_07291_));
 AND4_X1 _32323_ (.A1(_05696_),
    .A2(_05657_),
    .A3(_05525_),
    .A4(_05666_),
    .ZN(_07292_));
 AND3_X1 _32324_ (.A1(_05646_),
    .A2(_06242_),
    .A3(_05714_),
    .ZN(_07294_));
 AND2_X1 _32325_ (.A1(_05695_),
    .A2(_05631_),
    .ZN(_07295_));
 NOR4_X1 _32326_ (.A1(_07292_),
    .A2(_07294_),
    .A3(_07295_),
    .A4(_06696_),
    .ZN(_07296_));
 OAI21_X1 _32327_ (.A(_06711_),
    .B1(_06346_),
    .B2(_05575_),
    .ZN(_07297_));
 OAI211_X1 _32328_ (.A(_06711_),
    .B(_06285_),
    .C1(_05711_),
    .C2(_05611_),
    .ZN(_07298_));
 AND4_X1 _32329_ (.A1(_07291_),
    .A2(_07296_),
    .A3(_07297_),
    .A4(_07298_),
    .ZN(_07299_));
 AND3_X1 _32330_ (.A1(_05721_),
    .A2(_05589_),
    .A3(_05496_),
    .ZN(_07300_));
 AND2_X1 _32331_ (.A1(_05504_),
    .A2(_05498_),
    .ZN(_07301_));
 AND2_X1 _32332_ (.A1(_07301_),
    .A2(_05721_),
    .ZN(_07302_));
 AOI211_X1 _32333_ (.A(_07300_),
    .B(_07302_),
    .C1(_05703_),
    .C2(_05722_),
    .ZN(_07303_));
 OAI211_X1 _32334_ (.A(_06343_),
    .B(_05715_),
    .C1(_05713_),
    .C2(_05499_),
    .ZN(_07305_));
 OAI211_X1 _32335_ (.A(_05681_),
    .B(_06291_),
    .C1(_05711_),
    .C2(_05593_),
    .ZN(_07306_));
 OAI21_X1 _32336_ (.A(_06343_),
    .B1(_05633_),
    .B2(_05705_),
    .ZN(_07307_));
 OAI21_X1 _32337_ (.A(_06343_),
    .B1(_05557_),
    .B2(_06346_),
    .ZN(_07308_));
 AND4_X1 _32338_ (.A1(_07305_),
    .A2(_07306_),
    .A3(_07307_),
    .A4(_07308_),
    .ZN(_07309_));
 OAI21_X1 _32339_ (.A(_05722_),
    .B1(_06268_),
    .B2(_05543_),
    .ZN(_07310_));
 OAI211_X1 _32340_ (.A(_05722_),
    .B(_06291_),
    .C1(_05535_),
    .C2(_05572_),
    .ZN(_07311_));
 AND4_X1 _32341_ (.A1(_07303_),
    .A2(_07309_),
    .A3(_07310_),
    .A4(_07311_),
    .ZN(_07312_));
 NAND4_X1 _32342_ (.A1(_07277_),
    .A2(_07288_),
    .A3(_07299_),
    .A4(_07312_),
    .ZN(_07313_));
 AND3_X1 _32343_ (.A1(_05491_),
    .A2(_05496_),
    .A3(_05525_),
    .ZN(_07314_));
 AOI211_X1 _32344_ (.A(_07314_),
    .B(_05526_),
    .C1(_05491_),
    .C2(_05601_),
    .ZN(_07316_));
 AOI21_X1 _32345_ (.A(_05510_),
    .B1(_06244_),
    .B2(_06329_),
    .ZN(_07317_));
 AOI21_X1 _32346_ (.A(_07317_),
    .B1(_05491_),
    .B2(_05633_),
    .ZN(_07318_));
 OAI21_X1 _32347_ (.A(_05541_),
    .B1(_06268_),
    .B2(_05543_),
    .ZN(_07319_));
 NAND2_X1 _32348_ (.A1(_05530_),
    .A2(_05690_),
    .ZN(_07320_));
 AND2_X1 _32349_ (.A1(_07319_),
    .A2(_07320_),
    .ZN(_07321_));
 OAI21_X1 _32350_ (.A(_05541_),
    .B1(_05540_),
    .B2(_05557_),
    .ZN(_07322_));
 AND4_X1 _32351_ (.A1(_07316_),
    .A2(_07318_),
    .A3(_07321_),
    .A4(_07322_),
    .ZN(_07323_));
 AND2_X1 _32352_ (.A1(_05505_),
    .A2(_05590_),
    .ZN(_07324_));
 OAI21_X1 _32353_ (.A(_05626_),
    .B1(_05701_),
    .B2(_07324_),
    .ZN(_07325_));
 AND2_X1 _32354_ (.A1(_05534_),
    .A2(_05537_),
    .ZN(_07327_));
 OAI21_X1 _32355_ (.A(_05626_),
    .B1(_07327_),
    .B2(_05619_),
    .ZN(_07328_));
 AND2_X1 _32356_ (.A1(_06280_),
    .A2(_06723_),
    .ZN(_07329_));
 INV_X1 _32357_ (.A(_05655_),
    .ZN(_07330_));
 OAI21_X1 _32358_ (.A(_05606_),
    .B1(_07330_),
    .B2(_05612_),
    .ZN(_07331_));
 AND4_X1 _32359_ (.A1(_07325_),
    .A2(_07328_),
    .A3(_07329_),
    .A4(_07331_),
    .ZN(_07332_));
 OAI21_X1 _32360_ (.A(_05609_),
    .B1(_05624_),
    .B2(_05619_),
    .ZN(_07333_));
 NAND2_X1 _32361_ (.A1(_06266_),
    .A2(_05703_),
    .ZN(_07334_));
 NAND2_X1 _32362_ (.A1(_06266_),
    .A2(_05589_),
    .ZN(_07335_));
 AND4_X1 _32363_ (.A1(_06277_),
    .A2(_07333_),
    .A3(_07334_),
    .A4(_07335_),
    .ZN(_07336_));
 OAI21_X1 _32364_ (.A(_05583_),
    .B1(_06268_),
    .B2(_05543_),
    .ZN(_07338_));
 AND2_X1 _32365_ (.A1(_05492_),
    .A2(_05590_),
    .ZN(_07339_));
 OAI21_X1 _32366_ (.A(_05583_),
    .B1(_07301_),
    .B2(_07339_),
    .ZN(_07340_));
 AND4_X1 _32367_ (.A1(_06293_),
    .A2(_07336_),
    .A3(_07338_),
    .A4(_07340_),
    .ZN(_07341_));
 OAI21_X1 _32368_ (.A(_06251_),
    .B1(_05674_),
    .B2(_06267_),
    .ZN(_07342_));
 OAI211_X1 _32369_ (.A(_05554_),
    .B(_05623_),
    .C1(_05711_),
    .C2(_16721_),
    .ZN(_07343_));
 NAND2_X1 _32370_ (.A1(_05557_),
    .A2(_06251_),
    .ZN(_07344_));
 NAND2_X1 _32371_ (.A1(_05547_),
    .A2(_05628_),
    .ZN(_07345_));
 AND4_X1 _32372_ (.A1(_07342_),
    .A2(_07343_),
    .A3(_07344_),
    .A4(_07345_),
    .ZN(_07346_));
 NAND4_X1 _32373_ (.A1(_07323_),
    .A2(_07332_),
    .A3(_07341_),
    .A4(_07346_),
    .ZN(_07347_));
 NOR2_X2 _32374_ (.A1(_07313_),
    .A2(_07347_),
    .ZN(_07349_));
 XOR2_X1 _32375_ (.A(_07269_),
    .B(_07349_),
    .Z(_07350_));
 XNOR2_X1 _32376_ (.A(_07195_),
    .B(_07350_),
    .ZN(_07351_));
 XOR2_X1 _32377_ (.A(_07111_),
    .B(_07351_),
    .Z(_07352_));
 MUX2_X1 _32378_ (.A(_07022_),
    .B(_07352_),
    .S(_05069_),
    .Z(_00703_));
 MUX2_X1 _32379_ (.A(_16964_),
    .B(_16836_),
    .S(_03836_),
    .Z(_00761_));
 MUX2_X1 _32380_ (.A(_16965_),
    .B(_16837_),
    .S(_03836_),
    .Z(_00762_));
 XOR2_X1 _32381_ (.A(_17125_),
    .B(_16936_),
    .Z(_07353_));
 OAI211_X1 _32382_ (.A(_05562_),
    .B(_05525_),
    .C1(_05494_),
    .C2(_05611_),
    .ZN(_07354_));
 NAND2_X1 _32383_ (.A1(_06251_),
    .A2(_05558_),
    .ZN(_07355_));
 NAND4_X1 _32384_ (.A1(_05505_),
    .A2(_05499_),
    .A3(_05506_),
    .A4(_05561_),
    .ZN(_07357_));
 AND3_X1 _32385_ (.A1(_07354_),
    .A2(_07355_),
    .A3(_07357_),
    .ZN(_07358_));
 AOI21_X1 _32386_ (.A(_06245_),
    .B1(_06244_),
    .B2(_06329_),
    .ZN(_07359_));
 INV_X1 _32387_ (.A(_06267_),
    .ZN(_07360_));
 OAI21_X1 _32388_ (.A(_07320_),
    .B1(_06245_),
    .B2(_07360_),
    .ZN(_07361_));
 AND3_X1 _32389_ (.A1(_05618_),
    .A2(_06242_),
    .A3(_05506_),
    .ZN(_07362_));
 AND3_X1 _32390_ (.A1(_07301_),
    .A2(_06242_),
    .A3(_05506_),
    .ZN(_07363_));
 NOR4_X1 _32391_ (.A1(_07359_),
    .A2(_07361_),
    .A3(_07362_),
    .A4(_07363_),
    .ZN(_07364_));
 NAND2_X1 _32392_ (.A1(_06257_),
    .A2(_05490_),
    .ZN(_07365_));
 AND3_X1 _32393_ (.A1(_05490_),
    .A2(_05504_),
    .A3(_05572_),
    .ZN(_07366_));
 INV_X1 _32394_ (.A(_07366_),
    .ZN(_07368_));
 NAND3_X1 _32395_ (.A1(_05490_),
    .A2(_05524_),
    .A3(_05572_),
    .ZN(_07369_));
 AND4_X1 _32396_ (.A1(_07365_),
    .A2(_07368_),
    .A3(_06750_),
    .A4(_07369_),
    .ZN(_07370_));
 OAI21_X1 _32397_ (.A(_05554_),
    .B1(_05540_),
    .B2(_05493_),
    .ZN(_07371_));
 AND3_X1 _32398_ (.A1(_05551_),
    .A2(_06255_),
    .A3(_07371_),
    .ZN(_07372_));
 AND4_X1 _32399_ (.A1(_07358_),
    .A2(_07364_),
    .A3(_07370_),
    .A4(_07372_),
    .ZN(_07373_));
 AOI21_X1 _32400_ (.A(_06287_),
    .B1(_06675_),
    .B2(_06713_),
    .ZN(_07374_));
 NAND4_X1 _32401_ (.A1(_06273_),
    .A2(_05589_),
    .A3(_06309_),
    .A4(_05494_),
    .ZN(_07375_));
 OAI21_X1 _32402_ (.A(_07375_),
    .B1(_06287_),
    .B2(_05648_),
    .ZN(_07376_));
 AND2_X1 _32403_ (.A1(_06729_),
    .A2(_05625_),
    .ZN(_07377_));
 AND4_X1 _32404_ (.A1(_05715_),
    .A2(_06273_),
    .A3(_05572_),
    .A4(_05561_),
    .ZN(_07379_));
 NOR4_X1 _32405_ (.A1(_07374_),
    .A2(_07376_),
    .A3(_07377_),
    .A4(_07379_),
    .ZN(_07380_));
 AOI211_X1 _32406_ (.A(_06263_),
    .B(_05598_),
    .C1(_05515_),
    .C2(_05611_),
    .ZN(_07381_));
 AND2_X1 _32407_ (.A1(_06705_),
    .A2(_05606_),
    .ZN(_07382_));
 AND2_X1 _32408_ (.A1(_05606_),
    .A2(_05612_),
    .ZN(_07383_));
 AND2_X1 _32409_ (.A1(_05564_),
    .A2(_05597_),
    .ZN(_07384_));
 NOR4_X1 _32410_ (.A1(_07381_),
    .A2(_07382_),
    .A3(_07383_),
    .A4(_07384_),
    .ZN(_07385_));
 AND2_X1 _32411_ (.A1(_05609_),
    .A2(_05699_),
    .ZN(_07386_));
 AOI211_X1 _32412_ (.A(_05614_),
    .B(_07386_),
    .C1(_05609_),
    .C2(_05616_),
    .ZN(_07387_));
 AND4_X1 _32413_ (.A1(_05567_),
    .A2(_06273_),
    .A3(_05535_),
    .A4(_05488_),
    .ZN(_07388_));
 AND2_X1 _32414_ (.A1(_05674_),
    .A2(_05582_),
    .ZN(_07390_));
 AOI211_X1 _32415_ (.A(_07388_),
    .B(_07390_),
    .C1(_05564_),
    .C2(_05582_),
    .ZN(_07391_));
 OAI21_X1 _32416_ (.A(_05609_),
    .B1(_05605_),
    .B2(_05508_),
    .ZN(_07392_));
 AND4_X1 _32417_ (.A1(_06290_),
    .A2(_07387_),
    .A3(_07391_),
    .A4(_07392_),
    .ZN(_07393_));
 NAND4_X1 _32418_ (.A1(_07373_),
    .A2(_07380_),
    .A3(_07385_),
    .A4(_07393_),
    .ZN(_07394_));
 AND2_X1 _32419_ (.A1(_05672_),
    .A2(_05644_),
    .ZN(_07395_));
 AOI211_X1 _32420_ (.A(_07285_),
    .B(_07395_),
    .C1(_05646_),
    .C2(_05673_),
    .ZN(_07396_));
 OAI21_X1 _32421_ (.A(_05670_),
    .B1(_05699_),
    .B2(_05644_),
    .ZN(_07397_));
 OAI21_X1 _32422_ (.A(_05670_),
    .B1(_06697_),
    .B2(_05628_),
    .ZN(_07398_));
 AND4_X1 _32423_ (.A1(_05641_),
    .A2(_07396_),
    .A3(_07397_),
    .A4(_07398_),
    .ZN(_07399_));
 AOI21_X1 _32424_ (.A(_05718_),
    .B1(_06282_),
    .B2(_05585_),
    .ZN(_07401_));
 OAI21_X1 _32425_ (.A(_05695_),
    .B1(_06304_),
    .B2(_06346_),
    .ZN(_07402_));
 OAI21_X1 _32426_ (.A(_05695_),
    .B1(_05644_),
    .B2(_05616_),
    .ZN(_07403_));
 NAND3_X1 _32427_ (.A1(_05564_),
    .A2(_06242_),
    .A3(_05679_),
    .ZN(_07404_));
 NAND3_X1 _32428_ (.A1(_07402_),
    .A2(_07403_),
    .A3(_07404_),
    .ZN(_07405_));
 AOI211_X1 _32429_ (.A(_07401_),
    .B(_07405_),
    .C1(_06711_),
    .C2(_06715_),
    .ZN(_07406_));
 OAI211_X1 _32430_ (.A(_05721_),
    .B(_16722_),
    .C1(_16721_),
    .C2(_05499_),
    .ZN(_07407_));
 OAI21_X1 _32431_ (.A(_05681_),
    .B1(_05623_),
    .B2(_05516_),
    .ZN(_07408_));
 OAI21_X1 _32432_ (.A(_05681_),
    .B1(_05692_),
    .B2(_05704_),
    .ZN(_07409_));
 AND4_X1 _32433_ (.A1(_05725_),
    .A2(_07407_),
    .A3(_07408_),
    .A4(_07409_),
    .ZN(_07410_));
 OR2_X1 _32434_ (.A1(_05659_),
    .A2(_06307_),
    .ZN(_07412_));
 AOI21_X1 _32435_ (.A(_05649_),
    .B1(_06703_),
    .B2(_05565_),
    .ZN(_07413_));
 AOI21_X1 _32436_ (.A(_05652_),
    .B1(_05509_),
    .B2(_05655_),
    .ZN(_07414_));
 NAND2_X1 _32437_ (.A1(_05642_),
    .A2(_06271_),
    .ZN(_07415_));
 OAI21_X1 _32438_ (.A(_07415_),
    .B1(_05649_),
    .B2(_05509_),
    .ZN(_07416_));
 NOR4_X1 _32439_ (.A1(_07412_),
    .A2(_07413_),
    .A3(_07414_),
    .A4(_07416_),
    .ZN(_07417_));
 NAND4_X1 _32440_ (.A1(_07399_),
    .A2(_07406_),
    .A3(_07410_),
    .A4(_07417_),
    .ZN(_07418_));
 NOR2_X2 _32441_ (.A1(_07394_),
    .A2(_07418_),
    .ZN(_07419_));
 NAND2_X1 _32442_ (.A1(_06384_),
    .A2(_05312_),
    .ZN(_07420_));
 OR2_X1 _32443_ (.A1(_06374_),
    .A2(_05158_),
    .ZN(_07421_));
 AND2_X1 _32444_ (.A1(_06819_),
    .A2(_05163_),
    .ZN(_07423_));
 INV_X1 _32445_ (.A(_07423_),
    .ZN(_07424_));
 NAND3_X1 _32446_ (.A1(_05163_),
    .A2(_05138_),
    .A3(_05150_),
    .ZN(_07425_));
 AND4_X1 _32447_ (.A1(_07421_),
    .A2(_06803_),
    .A3(_07424_),
    .A4(_07425_),
    .ZN(_07426_));
 OAI211_X1 _32448_ (.A(_06384_),
    .B(_06410_),
    .C1(_05140_),
    .C2(_05166_),
    .ZN(_07427_));
 OAI21_X1 _32449_ (.A(_07243_),
    .B1(_06386_),
    .B2(_05195_),
    .ZN(_07428_));
 AOI21_X1 _32450_ (.A(_07428_),
    .B1(_05370_),
    .B2(_06384_),
    .ZN(_07429_));
 AND4_X1 _32451_ (.A1(_07420_),
    .A2(_07426_),
    .A3(_07427_),
    .A4(_07429_),
    .ZN(_07430_));
 OAI21_X1 _32452_ (.A(_05311_),
    .B1(_05384_),
    .B2(_05462_),
    .ZN(_07431_));
 OAI21_X1 _32453_ (.A(_05311_),
    .B1(_05252_),
    .B2(_05301_),
    .ZN(_07432_));
 OAI211_X1 _32454_ (.A(_05286_),
    .B(_05129_),
    .C1(_05207_),
    .C2(_05141_),
    .ZN(_07434_));
 NAND4_X1 _32455_ (.A1(_05286_),
    .A2(_05138_),
    .A3(_05129_),
    .A4(_05157_),
    .ZN(_07435_));
 AND4_X1 _32456_ (.A1(_07431_),
    .A2(_07432_),
    .A3(_07434_),
    .A4(_07435_),
    .ZN(_07436_));
 OAI21_X1 _32457_ (.A(_05297_),
    .B1(_05250_),
    .B2(_05446_),
    .ZN(_07437_));
 OAI211_X1 _32458_ (.A(_06394_),
    .B(_06767_),
    .C1(_05235_),
    .C2(_05142_),
    .ZN(_07438_));
 AND4_X1 _32459_ (.A1(_07234_),
    .A2(_07436_),
    .A3(_07437_),
    .A4(_07438_),
    .ZN(_07439_));
 INV_X1 _32460_ (.A(_05219_),
    .ZN(_07440_));
 OAI211_X1 _32461_ (.A(_05303_),
    .B(_05308_),
    .C1(_07263_),
    .C2(_07440_),
    .ZN(_07441_));
 AOI21_X1 _32462_ (.A(_07263_),
    .B1(_05454_),
    .B2(_06386_),
    .ZN(_07442_));
 AOI21_X1 _32463_ (.A(_05451_),
    .B1(_06408_),
    .B2(_05246_),
    .ZN(_07443_));
 NOR4_X1 _32464_ (.A1(_07441_),
    .A2(_07442_),
    .A3(_07443_),
    .A4(_06395_),
    .ZN(_07445_));
 OAI211_X1 _32465_ (.A(_05143_),
    .B(_05150_),
    .C1(_05140_),
    .C2(_05166_),
    .ZN(_07446_));
 OAI21_X1 _32466_ (.A(_05199_),
    .B1(_05183_),
    .B2(_05171_),
    .ZN(_07447_));
 OAI21_X1 _32467_ (.A(_05143_),
    .B1(_05370_),
    .B2(_05332_),
    .ZN(_07448_));
 OAI211_X1 _32468_ (.A(_05199_),
    .B(_05190_),
    .C1(_05200_),
    .C2(_05150_),
    .ZN(_07449_));
 AND4_X1 _32469_ (.A1(_07446_),
    .A2(_07447_),
    .A3(_07448_),
    .A4(_07449_),
    .ZN(_07450_));
 NAND4_X1 _32470_ (.A1(_07430_),
    .A2(_07439_),
    .A3(_07445_),
    .A4(_07450_),
    .ZN(_07451_));
 OAI21_X1 _32471_ (.A(_05262_),
    .B1(_05207_),
    .B2(_05142_),
    .ZN(_07452_));
 AND3_X1 _32472_ (.A1(_05372_),
    .A2(_05266_),
    .A3(_07452_),
    .ZN(_07453_));
 OAI21_X1 _32473_ (.A(_05244_),
    .B1(_05261_),
    .B2(_05177_),
    .ZN(_07454_));
 OAI21_X1 _32474_ (.A(_05244_),
    .B1(_05462_),
    .B2(_05256_),
    .ZN(_07456_));
 AND4_X1 _32475_ (.A1(_05461_),
    .A2(_07453_),
    .A3(_07454_),
    .A4(_07456_),
    .ZN(_07457_));
 INV_X1 _32476_ (.A(_06356_),
    .ZN(_07458_));
 OAI211_X1 _32477_ (.A(_07458_),
    .B(_07217_),
    .C1(_05400_),
    .C2(_05339_),
    .ZN(_07459_));
 NAND2_X1 _32478_ (.A1(_05334_),
    .A2(_05336_),
    .ZN(_07460_));
 AOI21_X1 _32479_ (.A(_05342_),
    .B1(_07440_),
    .B2(_05400_),
    .ZN(_07461_));
 NAND3_X1 _32480_ (.A1(_05204_),
    .A2(_05347_),
    .A3(_05190_),
    .ZN(_07462_));
 OAI21_X1 _32481_ (.A(_07462_),
    .B1(_05342_),
    .B2(_05378_),
    .ZN(_07463_));
 NOR4_X1 _32482_ (.A1(_07459_),
    .A2(_07460_),
    .A3(_07461_),
    .A4(_07463_),
    .ZN(_07464_));
 OAI211_X1 _32483_ (.A(_05220_),
    .B(_05168_),
    .C1(_05164_),
    .C2(_05166_),
    .ZN(_07465_));
 OAI21_X1 _32484_ (.A(_07465_),
    .B1(_07199_),
    .B2(_05239_),
    .ZN(_07467_));
 NAND2_X1 _32485_ (.A1(_05220_),
    .A2(_05284_),
    .ZN(_07468_));
 NAND3_X1 _32486_ (.A1(_05218_),
    .A2(_05469_),
    .A3(_07468_),
    .ZN(_07469_));
 AOI21_X1 _32487_ (.A(_05381_),
    .B1(_06408_),
    .B2(_05449_),
    .ZN(_07470_));
 NOR4_X1 _32488_ (.A1(_07467_),
    .A2(_07469_),
    .A3(_06783_),
    .A4(_07470_),
    .ZN(_07471_));
 AOI22_X1 _32489_ (.A1(_06368_),
    .A2(_05343_),
    .B1(_06372_),
    .B2(_05329_),
    .ZN(_07472_));
 OAI21_X1 _32490_ (.A(_05358_),
    .B1(_05362_),
    .B2(_06372_),
    .ZN(_07473_));
 OAI21_X1 _32491_ (.A(_05329_),
    .B1(_05446_),
    .B2(_05312_),
    .ZN(_07474_));
 AND4_X1 _32492_ (.A1(_06353_),
    .A2(_07472_),
    .A3(_07473_),
    .A4(_07474_),
    .ZN(_07475_));
 NAND4_X1 _32493_ (.A1(_07457_),
    .A2(_07464_),
    .A3(_07471_),
    .A4(_07475_),
    .ZN(_07476_));
 NOR2_X2 _32494_ (.A1(_07451_),
    .A2(_07476_),
    .ZN(_07478_));
 XOR2_X2 _32495_ (.A(_07419_),
    .B(_07478_),
    .Z(_07479_));
 XNOR2_X1 _32496_ (.A(_07479_),
    .B(_00993_),
    .ZN(_07480_));
 XOR2_X2 _32497_ (.A(_05484_),
    .B(_07269_),
    .Z(_07481_));
 XNOR2_X1 _32498_ (.A(_07480_),
    .B(_07481_),
    .ZN(_07482_));
 INV_X1 _32499_ (.A(_06565_),
    .ZN(_07483_));
 NAND2_X1 _32500_ (.A1(_05972_),
    .A2(_05807_),
    .ZN(_07484_));
 NAND2_X1 _32501_ (.A1(_07483_),
    .A2(_07484_),
    .ZN(_07485_));
 AND2_X1 _32502_ (.A1(_05974_),
    .A2(_05783_),
    .ZN(_07486_));
 NOR4_X1 _32503_ (.A1(_07485_),
    .A2(_07112_),
    .A3(_07486_),
    .A4(_06938_),
    .ZN(_07487_));
 NAND4_X1 _32504_ (.A1(_05948_),
    .A2(_05850_),
    .A3(_05802_),
    .A4(_05851_),
    .ZN(_07489_));
 OAI211_X1 _32505_ (.A(_05979_),
    .B(_05892_),
    .C1(_05780_),
    .C2(_06572_),
    .ZN(_07490_));
 AND2_X1 _32506_ (.A1(_05979_),
    .A2(_05878_),
    .ZN(_07491_));
 AND3_X1 _32507_ (.A1(_05979_),
    .A2(_05747_),
    .A3(_06660_),
    .ZN(_07492_));
 AOI211_X1 _32508_ (.A(_07491_),
    .B(_07492_),
    .C1(_06609_),
    .C2(_05979_),
    .ZN(_07493_));
 NAND4_X1 _32509_ (.A1(_07487_),
    .A2(_07489_),
    .A3(_07490_),
    .A4(_07493_),
    .ZN(_07494_));
 AND2_X1 _32510_ (.A1(_05938_),
    .A2(_05829_),
    .ZN(_07495_));
 INV_X1 _32511_ (.A(_07495_),
    .ZN(_07496_));
 NAND3_X1 _32512_ (.A1(_05939_),
    .A2(_05763_),
    .A3(_05892_),
    .ZN(_07497_));
 OAI211_X1 _32513_ (.A(_07496_),
    .B(_07497_),
    .C1(_06960_),
    .C2(_05960_),
    .ZN(_07498_));
 INV_X1 _32514_ (.A(_05931_),
    .ZN(_07500_));
 AOI21_X1 _32515_ (.A(_06960_),
    .B1(_07500_),
    .B2(_06987_),
    .ZN(_07501_));
 NOR4_X1 _32516_ (.A1(_07498_),
    .A2(_05944_),
    .A3(_06629_),
    .A4(_07501_),
    .ZN(_07502_));
 NAND3_X1 _32517_ (.A1(_05912_),
    .A2(_05779_),
    .A3(_05887_),
    .ZN(_07503_));
 OAI211_X1 _32518_ (.A(_05912_),
    .B(_05892_),
    .C1(_05767_),
    .C2(_05763_),
    .ZN(_07504_));
 OAI211_X1 _32519_ (.A(_05912_),
    .B(_05977_),
    .C1(_05850_),
    .C2(_06572_),
    .ZN(_07505_));
 OAI21_X1 _32520_ (.A(_05912_),
    .B1(_05937_),
    .B2(_05831_),
    .ZN(_07506_));
 AND4_X1 _32521_ (.A1(_07503_),
    .A2(_07504_),
    .A3(_07505_),
    .A4(_07506_),
    .ZN(_07507_));
 OAI211_X1 _32522_ (.A(_05900_),
    .B(_05851_),
    .C1(_05746_),
    .C2(_05887_),
    .ZN(_07508_));
 OAI211_X1 _32523_ (.A(_05900_),
    .B(_05892_),
    .C1(_05780_),
    .C2(_05781_),
    .ZN(_07509_));
 OAI211_X1 _32524_ (.A(_05900_),
    .B(_05833_),
    .C1(_05850_),
    .C2(_05781_),
    .ZN(_07511_));
 OAI21_X1 _32525_ (.A(_05900_),
    .B1(_06559_),
    .B2(_06609_),
    .ZN(_07512_));
 AND4_X1 _32526_ (.A1(_07508_),
    .A2(_07509_),
    .A3(_07511_),
    .A4(_07512_),
    .ZN(_07513_));
 OAI21_X1 _32527_ (.A(_06604_),
    .B1(_05765_),
    .B2(_05807_),
    .ZN(_07514_));
 NAND2_X1 _32528_ (.A1(_06604_),
    .A2(_06609_),
    .ZN(_07515_));
 NAND3_X1 _32529_ (.A1(_05864_),
    .A2(_05848_),
    .A3(_05906_),
    .ZN(_07516_));
 AND4_X1 _32530_ (.A1(_05933_),
    .A2(_07514_),
    .A3(_07515_),
    .A4(_07516_),
    .ZN(_07517_));
 NAND4_X1 _32531_ (.A1(_07502_),
    .A2(_07507_),
    .A3(_07513_),
    .A4(_07517_),
    .ZN(_07518_));
 AND2_X1 _32532_ (.A1(_06605_),
    .A2(_05958_),
    .ZN(_07519_));
 AND2_X1 _32533_ (.A1(_05958_),
    .A2(_05765_),
    .ZN(_07520_));
 AND2_X1 _32534_ (.A1(_05958_),
    .A2(_05866_),
    .ZN(_07522_));
 OR4_X1 _32535_ (.A1(_07141_),
    .A2(_07519_),
    .A3(_07520_),
    .A4(_07522_),
    .ZN(_07523_));
 AND2_X1 _32536_ (.A1(_05846_),
    .A2(_05952_),
    .ZN(_07524_));
 AND3_X1 _32537_ (.A1(_06618_),
    .A2(_05756_),
    .A3(_05948_),
    .ZN(_07525_));
 OR4_X1 _32538_ (.A1(_07524_),
    .A2(_06940_),
    .A3(_07132_),
    .A4(_07525_),
    .ZN(_07526_));
 NOR4_X1 _32539_ (.A1(_07494_),
    .A2(_07518_),
    .A3(_07523_),
    .A4(_07526_),
    .ZN(_07527_));
 AND2_X1 _32540_ (.A1(_05833_),
    .A2(_05780_),
    .ZN(_07528_));
 OAI21_X1 _32541_ (.A(_05809_),
    .B1(_05878_),
    .B2(_07528_),
    .ZN(_07529_));
 NOR3_X1 _32542_ (.A1(_06973_),
    .A2(_07159_),
    .A3(_06972_),
    .ZN(_07530_));
 OAI21_X1 _32543_ (.A(_05809_),
    .B1(_06608_),
    .B2(_07163_),
    .ZN(_07531_));
 NAND2_X1 _32544_ (.A1(_05827_),
    .A2(_05931_),
    .ZN(_07533_));
 NAND2_X1 _32545_ (.A1(_05827_),
    .A2(_05878_),
    .ZN(_07534_));
 AND4_X1 _32546_ (.A1(_05835_),
    .A2(_07533_),
    .A3(_07534_),
    .A4(_05838_),
    .ZN(_07535_));
 AND4_X1 _32547_ (.A1(_07529_),
    .A2(_07530_),
    .A3(_07531_),
    .A4(_07535_),
    .ZN(_07536_));
 OAI21_X1 _32548_ (.A(_05751_),
    .B1(_06608_),
    .B2(_05804_),
    .ZN(_07537_));
 AND2_X1 _32549_ (.A1(_05757_),
    .A2(_06568_),
    .ZN(_07538_));
 AND2_X1 _32550_ (.A1(_05771_),
    .A2(_05931_),
    .ZN(_07539_));
 AOI211_X1 _32551_ (.A(_07538_),
    .B(_07539_),
    .C1(_06559_),
    .C2(_05774_),
    .ZN(_07540_));
 AND3_X1 _32552_ (.A1(_05750_),
    .A2(_05767_),
    .A3(_05787_),
    .ZN(_07541_));
 AOI221_X4 _32553_ (.A(_07541_),
    .B1(_06559_),
    .B2(_05750_),
    .C1(_05887_),
    .C2(_07005_),
    .ZN(_07542_));
 NAND3_X1 _32554_ (.A1(_05771_),
    .A2(_05747_),
    .A3(_05851_),
    .ZN(_07544_));
 NAND2_X1 _32555_ (.A1(_05771_),
    .A2(_05811_),
    .ZN(_07545_));
 AND2_X1 _32556_ (.A1(_07544_),
    .A2(_07545_),
    .ZN(_07546_));
 AND4_X1 _32557_ (.A1(_07537_),
    .A2(_07540_),
    .A3(_07542_),
    .A4(_07546_),
    .ZN(_07547_));
 NAND2_X1 _32558_ (.A1(_05843_),
    .A2(_06618_),
    .ZN(_07548_));
 AND2_X1 _32559_ (.A1(_05842_),
    .A2(_05959_),
    .ZN(_07549_));
 INV_X1 _32560_ (.A(_07549_),
    .ZN(_07550_));
 NAND2_X1 _32561_ (.A1(_05842_),
    .A2(_05778_),
    .ZN(_07551_));
 OAI21_X1 _32562_ (.A(_05842_),
    .B1(_05866_),
    .B2(_05789_),
    .ZN(_07552_));
 AND4_X1 _32563_ (.A1(_07548_),
    .A2(_07550_),
    .A3(_07551_),
    .A4(_07552_),
    .ZN(_07553_));
 OAI211_X1 _32564_ (.A(_05861_),
    .B(_05851_),
    .C1(_05780_),
    .C2(_06572_),
    .ZN(_07555_));
 OAI21_X1 _32565_ (.A(_05861_),
    .B1(_05834_),
    .B2(_05913_),
    .ZN(_07556_));
 AND4_X1 _32566_ (.A1(_06983_),
    .A2(_07553_),
    .A3(_07555_),
    .A4(_07556_),
    .ZN(_07557_));
 INV_X1 _32567_ (.A(_05879_),
    .ZN(_07558_));
 OAI21_X1 _32568_ (.A(_06561_),
    .B1(_05864_),
    .B2(_06618_),
    .ZN(_07559_));
 NAND2_X1 _32569_ (.A1(_06559_),
    .A2(_05883_),
    .ZN(_07560_));
 NAND3_X1 _32570_ (.A1(_05744_),
    .A2(_05747_),
    .A3(_05886_),
    .ZN(_07561_));
 AND4_X1 _32571_ (.A1(_07558_),
    .A2(_07559_),
    .A3(_07560_),
    .A4(_07561_),
    .ZN(_07562_));
 AND4_X1 _32572_ (.A1(_07536_),
    .A2(_07547_),
    .A3(_07557_),
    .A4(_07562_),
    .ZN(_07563_));
 AND2_X2 _32573_ (.A1(_07527_),
    .A2(_07563_),
    .ZN(_07564_));
 XOR2_X2 _32574_ (.A(_07564_),
    .B(_05983_),
    .Z(_07566_));
 NAND2_X1 _32575_ (.A1(_06495_),
    .A2(_05997_),
    .ZN(_07567_));
 NAND2_X1 _32576_ (.A1(_06035_),
    .A2(_06860_),
    .ZN(_07568_));
 OR2_X1 _32577_ (.A1(_06871_),
    .A2(_06205_),
    .ZN(_07569_));
 OAI21_X1 _32578_ (.A(_06023_),
    .B1(_06086_),
    .B2(_06052_),
    .ZN(_07570_));
 AND4_X1 _32579_ (.A1(_07568_),
    .A2(_07569_),
    .A3(_06870_),
    .A4(_07570_),
    .ZN(_07571_));
 AOI21_X1 _32580_ (.A(_06867_),
    .B1(_06069_),
    .B2(_05997_),
    .ZN(_07572_));
 AND4_X1 _32581_ (.A1(_07567_),
    .A2(_07571_),
    .A3(_06476_),
    .A4(_07572_),
    .ZN(_07573_));
 AND3_X1 _32582_ (.A1(_06860_),
    .A2(_05994_),
    .A3(_06158_),
    .ZN(_07574_));
 AOI211_X1 _32583_ (.A(_07574_),
    .B(_06139_),
    .C1(_06146_),
    .C2(_06137_),
    .ZN(_07575_));
 OAI21_X1 _32584_ (.A(_06167_),
    .B1(_06101_),
    .B2(_06168_),
    .ZN(_07577_));
 NAND2_X1 _32585_ (.A1(_06167_),
    .A2(_06143_),
    .ZN(_07578_));
 AND2_X1 _32586_ (.A1(_07577_),
    .A2(_07578_),
    .ZN(_07579_));
 OAI21_X1 _32587_ (.A(_06167_),
    .B1(_06086_),
    .B2(_06482_),
    .ZN(_07580_));
 AND4_X1 _32588_ (.A1(_06503_),
    .A2(_07575_),
    .A3(_07579_),
    .A4(_07580_),
    .ZN(_07581_));
 NAND2_X1 _32589_ (.A1(_06153_),
    .A2(_06114_),
    .ZN(_07582_));
 NAND3_X1 _32590_ (.A1(_06153_),
    .A2(_06125_),
    .A3(_06124_),
    .ZN(_07583_));
 OAI211_X1 _32591_ (.A(_06153_),
    .B(_06059_),
    .C1(_06044_),
    .C2(_06065_),
    .ZN(_07584_));
 NAND4_X1 _32592_ (.A1(_06148_),
    .A2(_07582_),
    .A3(_07583_),
    .A4(_07584_),
    .ZN(_07585_));
 AND2_X1 _32593_ (.A1(_06844_),
    .A2(_06190_),
    .ZN(_07586_));
 AND2_X1 _32594_ (.A1(_06844_),
    .A2(_06007_),
    .ZN(_07588_));
 OAI211_X1 _32595_ (.A(_06158_),
    .B(_06183_),
    .C1(_06049_),
    .C2(_06889_),
    .ZN(_07589_));
 NAND2_X1 _32596_ (.A1(_06844_),
    .A2(_06091_),
    .ZN(_07590_));
 NAND3_X1 _32597_ (.A1(_07589_),
    .A2(_06846_),
    .A3(_07590_),
    .ZN(_07591_));
 NOR4_X1 _32598_ (.A1(_07585_),
    .A2(_07586_),
    .A3(_07588_),
    .A4(_07591_),
    .ZN(_07592_));
 OAI21_X1 _32599_ (.A(_06849_),
    .B1(_06069_),
    .B2(_06095_),
    .ZN(_07593_));
 AND3_X1 _32600_ (.A1(_06063_),
    .A2(_06198_),
    .A3(_06014_),
    .ZN(_07594_));
 AND3_X1 _32601_ (.A1(_07025_),
    .A2(_06007_),
    .A3(_06125_),
    .ZN(_07595_));
 AOI211_X1 _32602_ (.A(_07594_),
    .B(_07595_),
    .C1(_06049_),
    .C2(_07025_),
    .ZN(_07596_));
 OAI211_X1 _32603_ (.A(_06849_),
    .B(_05992_),
    .C1(_06007_),
    .C2(_06043_),
    .ZN(_07597_));
 OAI21_X1 _32604_ (.A(_06849_),
    .B1(_06049_),
    .B2(_06889_),
    .ZN(_07599_));
 AND4_X1 _32605_ (.A1(_07593_),
    .A2(_07596_),
    .A3(_07597_),
    .A4(_07599_),
    .ZN(_07600_));
 NAND4_X1 _32606_ (.A1(_07573_),
    .A2(_07581_),
    .A3(_07592_),
    .A4(_07600_),
    .ZN(_07601_));
 NAND2_X1 _32607_ (.A1(_06097_),
    .A2(_06146_),
    .ZN(_07602_));
 OAI21_X1 _32608_ (.A(_06097_),
    .B1(_06103_),
    .B2(_06143_),
    .ZN(_07603_));
 OAI211_X1 _32609_ (.A(_06097_),
    .B(_06014_),
    .C1(_06008_),
    .C2(_06009_),
    .ZN(_07604_));
 NAND4_X1 _32610_ (.A1(_06902_),
    .A2(_07602_),
    .A3(_07603_),
    .A4(_07604_),
    .ZN(_07605_));
 INV_X1 _32611_ (.A(_06484_),
    .ZN(_07606_));
 AOI21_X1 _32612_ (.A(_06117_),
    .B1(_07606_),
    .B2(_06851_),
    .ZN(_07607_));
 NOR3_X1 _32613_ (.A1(_07605_),
    .A2(_06910_),
    .A3(_07607_),
    .ZN(_07608_));
 INV_X1 _32614_ (.A(_06081_),
    .ZN(_07610_));
 OAI21_X1 _32615_ (.A(_06122_),
    .B1(_06495_),
    .B2(_06188_),
    .ZN(_07611_));
 OAI211_X1 _32616_ (.A(_06082_),
    .B(_16762_),
    .C1(_16761_),
    .C2(_06198_),
    .ZN(_07612_));
 OAI21_X1 _32617_ (.A(_06122_),
    .B1(_06099_),
    .B2(_06130_),
    .ZN(_07613_));
 AND4_X1 _32618_ (.A1(_07610_),
    .A2(_07611_),
    .A3(_07612_),
    .A4(_07613_),
    .ZN(_07614_));
 OAI21_X1 _32619_ (.A(_06197_),
    .B1(_06146_),
    .B2(_06860_),
    .ZN(_07615_));
 OAI21_X1 _32620_ (.A(_06197_),
    .B1(_06170_),
    .B2(_06889_),
    .ZN(_07616_));
 NAND4_X1 _32621_ (.A1(_06172_),
    .A2(_06014_),
    .A3(_06213_),
    .A4(_06008_),
    .ZN(_07617_));
 NAND3_X1 _32622_ (.A1(_07615_),
    .A2(_07616_),
    .A3(_07617_),
    .ZN(_07618_));
 AOI21_X1 _32623_ (.A(_06539_),
    .B1(_05989_),
    .B2(_06514_),
    .ZN(_07619_));
 NOR4_X1 _32624_ (.A1(_07618_),
    .A2(_06541_),
    .A3(_07619_),
    .A4(_06222_),
    .ZN(_07621_));
 INV_X1 _32625_ (.A(_06216_),
    .ZN(_07622_));
 OAI21_X1 _32626_ (.A(_07081_),
    .B1(_06101_),
    .B2(_06103_),
    .ZN(_07623_));
 OAI21_X1 _32627_ (.A(_06210_),
    .B1(_06200_),
    .B2(_06151_),
    .ZN(_07624_));
 OAI21_X1 _32628_ (.A(_07081_),
    .B1(_06522_),
    .B2(_06107_),
    .ZN(_07625_));
 AND4_X1 _32629_ (.A1(_07622_),
    .A2(_07623_),
    .A3(_07624_),
    .A4(_07625_),
    .ZN(_07626_));
 NAND4_X1 _32630_ (.A1(_07608_),
    .A2(_07614_),
    .A3(_07621_),
    .A4(_07626_),
    .ZN(_07627_));
 NOR2_X2 _32631_ (.A1(_07601_),
    .A2(_07627_),
    .ZN(_07628_));
 XOR2_X1 _32632_ (.A(_07566_),
    .B(_07628_),
    .Z(_07629_));
 XNOR2_X1 _32633_ (.A(_07482_),
    .B(_07629_),
    .ZN(_07630_));
 MUX2_X1 _32634_ (.A(_07353_),
    .B(_07630_),
    .S(_05069_),
    .Z(_00704_));
 XOR2_X1 _32635_ (.A(_17126_),
    .B(_16937_),
    .Z(_07632_));
 AND3_X1 _32636_ (.A1(_05491_),
    .A2(_05711_),
    .A3(_05525_),
    .ZN(_07633_));
 NAND2_X1 _32637_ (.A1(_06244_),
    .A2(_06247_),
    .ZN(_07634_));
 OAI21_X1 _32638_ (.A(_05626_),
    .B1(_07634_),
    .B2(_05701_),
    .ZN(_07635_));
 OAI211_X1 _32639_ (.A(_07635_),
    .B(_07365_),
    .C1(_06329_),
    .C2(_05510_),
    .ZN(_07636_));
 OAI211_X1 _32640_ (.A(_06255_),
    .B(_06737_),
    .C1(_05598_),
    .C2(_05568_),
    .ZN(_07637_));
 OR4_X1 _32641_ (.A1(_07633_),
    .A2(_07636_),
    .A3(_07314_),
    .A4(_07637_),
    .ZN(_07638_));
 AND2_X1 _32642_ (.A1(_05703_),
    .A2(_05491_),
    .ZN(_07639_));
 AOI22_X1 _32643_ (.A1(_05670_),
    .A2(_06731_),
    .B1(_05696_),
    .B2(_05633_),
    .ZN(_07640_));
 OAI221_X1 _32644_ (.A(_07640_),
    .B1(_05648_),
    .B2(_05510_),
    .C1(_07360_),
    .C2(_05663_),
    .ZN(_07642_));
 OAI22_X1 _32645_ (.A1(_05649_),
    .A2(_06675_),
    .B1(_06287_),
    .B2(_06249_),
    .ZN(_07643_));
 OR4_X1 _32646_ (.A1(_07639_),
    .A2(_07642_),
    .A3(_07383_),
    .A4(_07643_),
    .ZN(_07644_));
 AND2_X1 _32647_ (.A1(_05625_),
    .A2(_05646_),
    .ZN(_07645_));
 AND2_X1 _32648_ (.A1(_05645_),
    .A2(_05721_),
    .ZN(_07646_));
 OR3_X1 _32649_ (.A1(_07384_),
    .A2(_07645_),
    .A3(_07646_),
    .ZN(_07647_));
 AND3_X1 _32650_ (.A1(_05692_),
    .A2(_05596_),
    .A3(_06273_),
    .ZN(_07648_));
 INV_X1 _32651_ (.A(_05721_),
    .ZN(_07649_));
 INV_X1 _32652_ (.A(_07339_),
    .ZN(_07650_));
 OAI22_X1 _32653_ (.A1(_06287_),
    .A2(_06713_),
    .B1(_07649_),
    .B2(_07650_),
    .ZN(_07651_));
 OR4_X1 _32654_ (.A1(_07275_),
    .A2(_07647_),
    .A3(_07648_),
    .A4(_07651_),
    .ZN(_07653_));
 NOR2_X1 _32655_ (.A1(_05658_),
    .A2(_05498_),
    .ZN(_07654_));
 NAND2_X1 _32656_ (.A1(_07654_),
    .A2(_05530_),
    .ZN(_07655_));
 NAND3_X1 _32657_ (.A1(_05575_),
    .A2(_06309_),
    .A3(_06312_),
    .ZN(_07656_));
 OAI211_X1 _32658_ (.A(_07655_),
    .B(_07656_),
    .C1(_06324_),
    .C2(_05585_),
    .ZN(_07657_));
 NOR4_X1 _32659_ (.A1(_07638_),
    .A2(_07644_),
    .A3(_07653_),
    .A4(_07657_),
    .ZN(_07658_));
 NAND4_X1 _32660_ (.A1(_06271_),
    .A2(_05666_),
    .A3(_05716_),
    .A4(_05638_),
    .ZN(_07659_));
 NAND4_X1 _32661_ (.A1(_05638_),
    .A2(_05505_),
    .A3(_05499_),
    .A4(_05488_),
    .ZN(_07660_));
 OAI211_X1 _32662_ (.A(_07659_),
    .B(_07660_),
    .C1(_05509_),
    .C2(_05652_),
    .ZN(_07661_));
 AOI221_X4 _32663_ (.A(_07661_),
    .B1(_05619_),
    .B2(_05651_),
    .C1(_05583_),
    .C2(_05594_),
    .ZN(_07662_));
 OAI21_X1 _32664_ (.A(_06343_),
    .B1(_07634_),
    .B2(_05587_),
    .ZN(_07664_));
 OAI21_X1 _32665_ (.A(_06266_),
    .B1(_05564_),
    .B2(_05690_),
    .ZN(_07665_));
 OAI21_X1 _32666_ (.A(_06266_),
    .B1(_06731_),
    .B2(_05703_),
    .ZN(_07666_));
 AND3_X1 _32667_ (.A1(_07665_),
    .A2(_07666_),
    .A3(_05620_),
    .ZN(_07667_));
 OR2_X1 _32668_ (.A1(_05701_),
    .A2(_06731_),
    .ZN(_07668_));
 NAND2_X1 _32669_ (.A1(_06244_),
    .A2(_05509_),
    .ZN(_07669_));
 OAI21_X1 _32670_ (.A(_05541_),
    .B1(_07668_),
    .B2(_07669_),
    .ZN(_07670_));
 NAND4_X1 _32671_ (.A1(_07662_),
    .A2(_07664_),
    .A3(_07667_),
    .A4(_07670_),
    .ZN(_07671_));
 AOI21_X1 _32672_ (.A(_05548_),
    .B1(_06249_),
    .B2(_05509_),
    .ZN(_07672_));
 AOI211_X1 _32673_ (.A(_05733_),
    .B(_07672_),
    .C1(_05554_),
    .C2(_07339_),
    .ZN(_07673_));
 OAI21_X1 _32674_ (.A(_06711_),
    .B1(_05701_),
    .B2(_07324_),
    .ZN(_07675_));
 OAI21_X1 _32675_ (.A(_06711_),
    .B1(_05543_),
    .B2(_05616_),
    .ZN(_07676_));
 NAND4_X1 _32676_ (.A1(_06711_),
    .A2(_06291_),
    .A3(_05537_),
    .A4(_05532_),
    .ZN(_07677_));
 AND3_X1 _32677_ (.A1(_07675_),
    .A2(_07676_),
    .A3(_07677_),
    .ZN(_07678_));
 AND2_X1 _32678_ (.A1(_07669_),
    .A2(_05662_),
    .ZN(_07679_));
 AND4_X1 _32679_ (.A1(_05611_),
    .A2(_06291_),
    .A3(_06273_),
    .A4(_05716_),
    .ZN(_07680_));
 AND4_X1 _32680_ (.A1(_05713_),
    .A2(_06273_),
    .A3(_05715_),
    .A4(_05716_),
    .ZN(_07681_));
 NOR3_X1 _32681_ (.A1(_07679_),
    .A2(_07680_),
    .A3(_07681_),
    .ZN(_07682_));
 AND2_X1 _32682_ (.A1(_05633_),
    .A2(_06251_),
    .ZN(_07683_));
 INV_X1 _32683_ (.A(_07683_),
    .ZN(_07684_));
 OAI21_X1 _32684_ (.A(_06251_),
    .B1(_06346_),
    .B2(_05575_),
    .ZN(_07686_));
 NAND4_X1 _32685_ (.A1(_05713_),
    .A2(_05715_),
    .A3(_06309_),
    .A4(_05506_),
    .ZN(_07687_));
 AND3_X1 _32686_ (.A1(_07684_),
    .A2(_07686_),
    .A3(_07687_),
    .ZN(_07688_));
 NAND4_X1 _32687_ (.A1(_07673_),
    .A2(_07678_),
    .A3(_07682_),
    .A4(_07688_),
    .ZN(_07689_));
 AND2_X1 _32688_ (.A1(_05642_),
    .A2(_06268_),
    .ZN(_07690_));
 OR4_X1 _32689_ (.A1(_05668_),
    .A2(_07690_),
    .A3(_07366_),
    .A4(_07362_),
    .ZN(_07691_));
 AOI22_X1 _32690_ (.A1(_05713_),
    .A2(_06291_),
    .B1(_06285_),
    .B2(_05711_),
    .ZN(_07692_));
 AOI21_X1 _32691_ (.A(_06324_),
    .B1(_06261_),
    .B2(_07692_),
    .ZN(_07693_));
 NAND2_X1 _32692_ (.A1(_05673_),
    .A2(_05644_),
    .ZN(_07694_));
 NAND4_X1 _32693_ (.A1(_06312_),
    .A2(_05713_),
    .A3(_05525_),
    .A4(_05596_),
    .ZN(_07695_));
 OAI211_X1 _32694_ (.A(_07694_),
    .B(_07695_),
    .C1(_06319_),
    .C2(_05585_),
    .ZN(_07697_));
 AOI21_X1 _32695_ (.A(_06319_),
    .B1(_05648_),
    .B2(_05509_),
    .ZN(_07698_));
 AOI21_X1 _32696_ (.A(_07649_),
    .B1(_06341_),
    .B2(_05658_),
    .ZN(_07699_));
 OR4_X1 _32697_ (.A1(_07693_),
    .A2(_07697_),
    .A3(_07698_),
    .A4(_07699_),
    .ZN(_07700_));
 NOR4_X1 _32698_ (.A1(_07671_),
    .A2(_07689_),
    .A3(_07691_),
    .A4(_07700_),
    .ZN(_07701_));
 AND2_X2 _32699_ (.A1(_07658_),
    .A2(_07701_),
    .ZN(_07702_));
 OAI21_X1 _32700_ (.A(_07255_),
    .B1(_05432_),
    .B2(_05249_),
    .ZN(_07703_));
 AOI221_X4 _32701_ (.A(_07703_),
    .B1(_05213_),
    .B2(_05143_),
    .C1(_05389_),
    .C2(_05263_),
    .ZN(_07704_));
 AOI22_X1 _32702_ (.A1(_05384_),
    .A2(_05263_),
    .B1(_05332_),
    .B2(_05175_),
    .ZN(_07705_));
 AND4_X1 _32703_ (.A1(_07421_),
    .A2(_07704_),
    .A3(_07420_),
    .A4(_07705_),
    .ZN(_07706_));
 OAI21_X1 _32704_ (.A(_06384_),
    .B1(_06360_),
    .B2(_06372_),
    .ZN(_07708_));
 OAI21_X1 _32705_ (.A(_06354_),
    .B1(_05213_),
    .B2(_05284_),
    .ZN(_07709_));
 OAI21_X1 _32706_ (.A(_06354_),
    .B1(_06372_),
    .B2(_05332_),
    .ZN(_07710_));
 NAND4_X1 _32707_ (.A1(_06767_),
    .A2(_05146_),
    .A3(_06410_),
    .A4(_05438_),
    .ZN(_07711_));
 AND3_X1 _32708_ (.A1(_07709_),
    .A2(_07710_),
    .A3(_07711_),
    .ZN(_07712_));
 NAND2_X1 _32709_ (.A1(_05389_),
    .A2(_05347_),
    .ZN(_07713_));
 NAND2_X1 _32710_ (.A1(_05311_),
    .A2(_05261_),
    .ZN(_07714_));
 AND4_X1 _32711_ (.A1(_07713_),
    .A2(_07714_),
    .A3(_05469_),
    .A4(_07242_),
    .ZN(_07715_));
 AND4_X1 _32712_ (.A1(_05319_),
    .A2(_07708_),
    .A3(_07712_),
    .A4(_07715_),
    .ZN(_07716_));
 NOR2_X1 _32713_ (.A1(_06367_),
    .A2(_06373_),
    .ZN(_07717_));
 OAI21_X1 _32714_ (.A(_05263_),
    .B1(_05252_),
    .B2(_05414_),
    .ZN(_07719_));
 AND4_X1 _32715_ (.A1(_05386_),
    .A2(_05367_),
    .A3(_07719_),
    .A4(_05264_),
    .ZN(_07720_));
 NAND3_X1 _32716_ (.A1(_05297_),
    .A2(_05155_),
    .A3(_05200_),
    .ZN(_07721_));
 NAND3_X1 _32717_ (.A1(_05177_),
    .A2(_05215_),
    .A3(_05267_),
    .ZN(_07722_));
 AND3_X1 _32718_ (.A1(_07721_),
    .A2(_06827_),
    .A3(_07722_),
    .ZN(_07723_));
 AND4_X1 _32719_ (.A1(_07717_),
    .A2(_07720_),
    .A3(_06830_),
    .A4(_07723_),
    .ZN(_07724_));
 NAND3_X1 _32720_ (.A1(_05194_),
    .A2(_07239_),
    .A3(_05378_),
    .ZN(_07725_));
 OAI21_X1 _32721_ (.A(_05380_),
    .B1(_07725_),
    .B2(_05200_),
    .ZN(_07726_));
 OAI21_X1 _32722_ (.A(_05441_),
    .B1(_05446_),
    .B2(_05252_),
    .ZN(_07727_));
 OAI21_X1 _32723_ (.A(_05441_),
    .B1(_06819_),
    .B2(_06372_),
    .ZN(_07728_));
 AND3_X1 _32724_ (.A1(_05305_),
    .A2(_07727_),
    .A3(_07728_),
    .ZN(_07730_));
 OAI21_X1 _32725_ (.A(_05358_),
    .B1(_05458_),
    .B2(_05204_),
    .ZN(_07731_));
 OAI21_X1 _32726_ (.A(_05244_),
    .B1(_05235_),
    .B2(_05316_),
    .ZN(_07732_));
 NAND4_X1 _32727_ (.A1(_06767_),
    .A2(_05138_),
    .A3(_06410_),
    .A4(_05267_),
    .ZN(_07733_));
 AND3_X1 _32728_ (.A1(_07732_),
    .A2(_05460_),
    .A3(_07733_),
    .ZN(_07734_));
 AND4_X1 _32729_ (.A1(_07726_),
    .A2(_07730_),
    .A3(_07731_),
    .A4(_07734_),
    .ZN(_07735_));
 NAND4_X1 _32730_ (.A1(_07706_),
    .A2(_07716_),
    .A3(_07724_),
    .A4(_07735_),
    .ZN(_07736_));
 AND2_X1 _32731_ (.A1(_05311_),
    .A2(_05301_),
    .ZN(_07737_));
 AND2_X1 _32732_ (.A1(_05347_),
    .A2(_05142_),
    .ZN(_07738_));
 OR4_X1 _32733_ (.A1(_05424_),
    .A2(_07737_),
    .A3(_05349_),
    .A4(_07738_),
    .ZN(_07739_));
 OAI21_X1 _32734_ (.A(_05199_),
    .B1(_06372_),
    .B2(_05414_),
    .ZN(_07741_));
 NAND3_X1 _32735_ (.A1(_07741_),
    .A2(_07468_),
    .A3(_07234_),
    .ZN(_07742_));
 OAI221_X1 _32736_ (.A(_05231_),
    .B1(_07199_),
    .B2(_05154_),
    .C1(_05292_),
    .C2(_05257_),
    .ZN(_07743_));
 NOR4_X1 _32737_ (.A1(_07739_),
    .A2(_05476_),
    .A3(_07742_),
    .A4(_07743_),
    .ZN(_07744_));
 OAI21_X1 _32738_ (.A(_05143_),
    .B1(_05316_),
    .B2(_05142_),
    .ZN(_07745_));
 AND2_X1 _32739_ (.A1(_05358_),
    .A2(_05312_),
    .ZN(_07746_));
 AOI21_X1 _32740_ (.A(_07746_),
    .B1(_05347_),
    .B2(_06819_),
    .ZN(_07747_));
 AOI21_X1 _32741_ (.A(_07423_),
    .B1(_05446_),
    .B2(_05297_),
    .ZN(_07748_));
 OAI21_X1 _32742_ (.A(_05281_),
    .B1(_05213_),
    .B2(_05320_),
    .ZN(_07749_));
 AND4_X1 _32743_ (.A1(_07745_),
    .A2(_07747_),
    .A3(_07748_),
    .A4(_07749_),
    .ZN(_07750_));
 AOI21_X1 _32744_ (.A(_05419_),
    .B1(_05430_),
    .B2(_05329_),
    .ZN(_07752_));
 OAI21_X1 _32745_ (.A(_06390_),
    .B1(_05199_),
    .B2(_05175_),
    .ZN(_07753_));
 AND3_X1 _32746_ (.A1(_07753_),
    .A2(_05287_),
    .A3(_05282_),
    .ZN(_07754_));
 NAND4_X1 _32747_ (.A1(_07744_),
    .A2(_07750_),
    .A3(_07752_),
    .A4(_07754_),
    .ZN(_07755_));
 NOR2_X2 _32748_ (.A1(_07736_),
    .A2(_07755_),
    .ZN(_07756_));
 XNOR2_X1 _32749_ (.A(_07702_),
    .B(_07756_),
    .ZN(_07757_));
 AND2_X1 _32750_ (.A1(_06210_),
    .A2(_06076_),
    .ZN(_07758_));
 AND2_X1 _32751_ (.A1(_06146_),
    .A2(_06210_),
    .ZN(_07759_));
 AND2_X1 _32752_ (.A1(_06209_),
    .A2(_06103_),
    .ZN(_07760_));
 AND2_X1 _32753_ (.A1(_06209_),
    .A2(_06190_),
    .ZN(_07761_));
 NOR4_X1 _32754_ (.A1(_07758_),
    .A2(_07759_),
    .A3(_07760_),
    .A4(_07761_),
    .ZN(_07763_));
 AOI21_X1 _32755_ (.A(_06206_),
    .B1(_06872_),
    .B2(_06514_),
    .ZN(_07764_));
 AND2_X1 _32756_ (.A1(_06086_),
    .A2(_06202_),
    .ZN(_07765_));
 NOR4_X1 _32757_ (.A1(_07764_),
    .A2(_07765_),
    .A3(_07080_),
    .A4(_06218_),
    .ZN(_07766_));
 OAI221_X1 _32758_ (.A(_06210_),
    .B1(_06032_),
    .B2(_06150_),
    .C1(_06014_),
    .C2(_06059_),
    .ZN(_07767_));
 NAND2_X1 _32759_ (.A1(_06151_),
    .A2(_07081_),
    .ZN(_07768_));
 AND2_X1 _32760_ (.A1(_06203_),
    .A2(_07768_),
    .ZN(_07769_));
 AND4_X1 _32761_ (.A1(_07763_),
    .A2(_07766_),
    .A3(_07767_),
    .A4(_07769_),
    .ZN(_07770_));
 NAND2_X1 _32762_ (.A1(_06224_),
    .A2(_06860_),
    .ZN(_07771_));
 OAI21_X1 _32763_ (.A(_06224_),
    .B1(_06510_),
    .B2(_06055_),
    .ZN(_07772_));
 OAI21_X1 _32764_ (.A(_06197_),
    .B1(_06128_),
    .B2(_06190_),
    .ZN(_07774_));
 AND4_X1 _32765_ (.A1(_07771_),
    .A2(_07036_),
    .A3(_07772_),
    .A4(_07774_),
    .ZN(_07775_));
 INV_X1 _32766_ (.A(_06096_),
    .ZN(_07776_));
 OAI21_X1 _32767_ (.A(_07776_),
    .B1(_06464_),
    .B2(_06098_),
    .ZN(_07777_));
 NAND4_X1 _32768_ (.A1(_06111_),
    .A2(_06007_),
    .A3(_05992_),
    .A4(_05987_),
    .ZN(_07778_));
 OAI211_X1 _32769_ (.A(_07778_),
    .B(_06914_),
    .C1(_06851_),
    .C2(_06117_),
    .ZN(_07779_));
 NAND2_X1 _32770_ (.A1(_06097_),
    .A2(_06000_),
    .ZN(_07780_));
 OAI211_X1 _32771_ (.A(_07780_),
    .B(_07602_),
    .C1(_06464_),
    .C2(_06851_),
    .ZN(_07781_));
 INV_X1 _32772_ (.A(_06106_),
    .ZN(_07782_));
 INV_X1 _32773_ (.A(_07070_),
    .ZN(_07783_));
 AOI21_X1 _32774_ (.A(_06117_),
    .B1(_07782_),
    .B2(_07783_),
    .ZN(_07785_));
 NOR4_X1 _32775_ (.A1(_07777_),
    .A2(_07779_),
    .A3(_07781_),
    .A4(_07785_),
    .ZN(_07786_));
 NAND2_X1 _32776_ (.A1(_06076_),
    .A2(_06082_),
    .ZN(_07787_));
 AND2_X1 _32777_ (.A1(_06151_),
    .A2(_06078_),
    .ZN(_07788_));
 INV_X1 _32778_ (.A(_07788_),
    .ZN(_07789_));
 NAND3_X1 _32779_ (.A1(_06450_),
    .A2(_07787_),
    .A3(_07789_),
    .ZN(_07790_));
 OAI21_X1 _32780_ (.A(_06122_),
    .B1(_06086_),
    .B2(_06095_),
    .ZN(_07791_));
 NAND2_X1 _32781_ (.A1(_06080_),
    .A2(_06122_),
    .ZN(_07792_));
 OAI211_X1 _32782_ (.A(_07791_),
    .B(_07792_),
    .C1(_06851_),
    .C2(_06120_),
    .ZN(_07793_));
 AND2_X1 _32783_ (.A1(_06082_),
    .A2(_07090_),
    .ZN(_07794_));
 AND3_X1 _32784_ (.A1(_06082_),
    .A2(_06032_),
    .A3(_06014_),
    .ZN(_07796_));
 NOR4_X1 _32785_ (.A1(_07790_),
    .A2(_07793_),
    .A3(_07794_),
    .A4(_07796_),
    .ZN(_07797_));
 NAND4_X1 _32786_ (.A1(_07770_),
    .A2(_07775_),
    .A3(_07786_),
    .A4(_07797_),
    .ZN(_07798_));
 AND2_X1 _32787_ (.A1(_06035_),
    .A2(_06069_),
    .ZN(_07799_));
 AOI211_X1 _32788_ (.A(_06483_),
    .B(_07799_),
    .C1(_06923_),
    .C2(_06035_),
    .ZN(_07800_));
 AND4_X1 _32789_ (.A1(_07567_),
    .A2(_06475_),
    .A3(_06476_),
    .A4(_06477_),
    .ZN(_07801_));
 OAI221_X1 _32790_ (.A(_05997_),
    .B1(_06008_),
    .B2(_06065_),
    .C1(_06014_),
    .C2(_06059_),
    .ZN(_07802_));
 OAI21_X1 _32791_ (.A(_06035_),
    .B1(_07026_),
    .B2(_06860_),
    .ZN(_07803_));
 NAND4_X1 _32792_ (.A1(_07800_),
    .A2(_07801_),
    .A3(_07802_),
    .A4(_07803_),
    .ZN(_07804_));
 AND2_X1 _32793_ (.A1(_06889_),
    .A2(_07025_),
    .ZN(_07805_));
 AND2_X1 _32794_ (.A1(_06095_),
    .A2(_07025_),
    .ZN(_07807_));
 AOI211_X1 _32795_ (.A(_07805_),
    .B(_07807_),
    .C1(_06049_),
    .C2(_07025_),
    .ZN(_07808_));
 NAND2_X1 _32796_ (.A1(_06103_),
    .A2(_07025_),
    .ZN(_07809_));
 OAI21_X1 _32797_ (.A(_06849_),
    .B1(_07090_),
    .B2(_06014_),
    .ZN(_07810_));
 OAI21_X1 _32798_ (.A(_06849_),
    .B1(_06019_),
    .B2(_06177_),
    .ZN(_07811_));
 NAND4_X1 _32799_ (.A1(_07808_),
    .A2(_07809_),
    .A3(_07810_),
    .A4(_07811_),
    .ZN(_07812_));
 OAI21_X1 _32800_ (.A(_07582_),
    .B1(_06161_),
    .B2(_06885_),
    .ZN(_07813_));
 NOR3_X1 _32801_ (.A1(_07813_),
    .A2(_06147_),
    .A3(_06513_),
    .ZN(_07814_));
 AOI21_X1 _32802_ (.A(_06140_),
    .B1(_06459_),
    .B2(_06540_),
    .ZN(_07815_));
 NOR2_X1 _32803_ (.A1(_07815_),
    .A2(_06142_),
    .ZN(_07816_));
 OAI21_X1 _32804_ (.A(_06018_),
    .B1(_06198_),
    .B2(_06025_),
    .ZN(_07818_));
 OAI21_X1 _32805_ (.A(_06167_),
    .B1(_07818_),
    .B2(_06860_),
    .ZN(_07819_));
 OAI21_X1 _32806_ (.A(_06844_),
    .B1(_06076_),
    .B2(_06168_),
    .ZN(_07820_));
 AND4_X1 _32807_ (.A1(_06181_),
    .A2(_07820_),
    .A3(_06184_),
    .A4(_06846_),
    .ZN(_07821_));
 NAND4_X1 _32808_ (.A1(_07814_),
    .A2(_07816_),
    .A3(_07819_),
    .A4(_07821_),
    .ZN(_07822_));
 NOR4_X1 _32809_ (.A1(_07798_),
    .A2(_07804_),
    .A3(_07812_),
    .A4(_07822_),
    .ZN(_07823_));
 INV_X1 _32810_ (.A(_06232_),
    .ZN(_07824_));
 NAND2_X2 _32811_ (.A1(_07823_),
    .A2(_07824_),
    .ZN(_07825_));
 XNOR2_X1 _32812_ (.A(_07825_),
    .B(_00994_),
    .ZN(_07826_));
 XOR2_X1 _32813_ (.A(_07757_),
    .B(_07826_),
    .Z(_07827_));
 AOI211_X1 _32814_ (.A(_07495_),
    .B(_07151_),
    .C1(_06977_),
    .C2(_05939_),
    .ZN(_07829_));
 AND2_X1 _32815_ (.A1(_06604_),
    .A2(_05829_),
    .ZN(_07830_));
 NOR3_X1 _32816_ (.A1(_05926_),
    .A2(_05927_),
    .A3(_07830_),
    .ZN(_07831_));
 OAI211_X1 _32817_ (.A(_06604_),
    .B(_05977_),
    .C1(_05850_),
    .C2(_06572_),
    .ZN(_07832_));
 AND4_X1 _32818_ (.A1(_07515_),
    .A2(_07829_),
    .A3(_07831_),
    .A4(_07832_),
    .ZN(_07833_));
 AND2_X1 _32819_ (.A1(_05765_),
    .A2(_05912_),
    .ZN(_07834_));
 INV_X1 _32820_ (.A(_07834_),
    .ZN(_07835_));
 OAI21_X1 _32821_ (.A(_05900_),
    .B1(_06575_),
    .B2(_06618_),
    .ZN(_07836_));
 OAI211_X1 _32822_ (.A(_05912_),
    .B(_16802_),
    .C1(_16801_),
    .C2(_05746_),
    .ZN(_07837_));
 OAI21_X1 _32823_ (.A(_05900_),
    .B1(_05789_),
    .B2(_05867_),
    .ZN(_07838_));
 AND4_X1 _32824_ (.A1(_07835_),
    .A2(_07836_),
    .A3(_07837_),
    .A4(_07838_),
    .ZN(_07840_));
 NAND2_X1 _32825_ (.A1(_06940_),
    .A2(_06662_),
    .ZN(_07841_));
 INV_X1 _32826_ (.A(_07522_),
    .ZN(_07842_));
 AND4_X1 _32827_ (.A1(_06614_),
    .A2(_07842_),
    .A3(_06932_),
    .A4(_06933_),
    .ZN(_07843_));
 OAI21_X1 _32828_ (.A(_05952_),
    .B1(_05857_),
    .B2(_07163_),
    .ZN(_07844_));
 NAND4_X1 _32829_ (.A1(_05848_),
    .A2(_05948_),
    .A3(_05977_),
    .A4(_06572_),
    .ZN(_07845_));
 AND4_X1 _32830_ (.A1(_07841_),
    .A2(_07843_),
    .A3(_07844_),
    .A4(_07845_),
    .ZN(_07846_));
 OAI21_X1 _32831_ (.A(_05974_),
    .B1(_05773_),
    .B2(_05864_),
    .ZN(_07847_));
 NAND4_X1 _32832_ (.A1(_07847_),
    .A2(_06612_),
    .A3(_06613_),
    .A4(_07484_),
    .ZN(_07848_));
 AOI21_X1 _32833_ (.A(_06591_),
    .B1(_06647_),
    .B2(_06997_),
    .ZN(_07849_));
 AND2_X1 _32834_ (.A1(_05846_),
    .A2(_05979_),
    .ZN(_07851_));
 NOR4_X1 _32835_ (.A1(_07848_),
    .A2(_07849_),
    .A3(_07851_),
    .A4(_07491_),
    .ZN(_07852_));
 NAND4_X1 _32836_ (.A1(_07833_),
    .A2(_07840_),
    .A3(_07846_),
    .A4(_07852_),
    .ZN(_07853_));
 INV_X1 _32837_ (.A(_06623_),
    .ZN(_07854_));
 NAND2_X1 _32838_ (.A1(_05843_),
    .A2(_05855_),
    .ZN(_07855_));
 NAND2_X1 _32839_ (.A1(_05843_),
    .A2(_05829_),
    .ZN(_07856_));
 AND3_X1 _32840_ (.A1(_07854_),
    .A2(_07855_),
    .A3(_07856_),
    .ZN(_07857_));
 OAI21_X1 _32841_ (.A(_05861_),
    .B1(_06977_),
    .B2(_07163_),
    .ZN(_07858_));
 OAI21_X1 _32842_ (.A(_05843_),
    .B1(_05969_),
    .B2(_05866_),
    .ZN(_07859_));
 AND4_X1 _32843_ (.A1(_06981_),
    .A2(_07857_),
    .A3(_07858_),
    .A4(_07859_),
    .ZN(_07860_));
 OAI21_X1 _32844_ (.A(_05828_),
    .B1(_05963_),
    .B2(_05857_),
    .ZN(_07862_));
 OAI211_X1 _32845_ (.A(_05828_),
    .B(_05779_),
    .C1(_05780_),
    .C2(_05781_),
    .ZN(_07863_));
 NAND4_X1 _32846_ (.A1(_07862_),
    .A2(_05835_),
    .A3(_07533_),
    .A4(_07863_),
    .ZN(_07864_));
 AND2_X1 _32847_ (.A1(_05809_),
    .A2(_05779_),
    .ZN(_07865_));
 OAI22_X1 _32848_ (.A1(_05740_),
    .A2(_05813_),
    .B1(_06571_),
    .B2(_06572_),
    .ZN(_07866_));
 NOR4_X1 _32849_ (.A1(_07864_),
    .A2(_05820_),
    .A3(_07865_),
    .A4(_07866_),
    .ZN(_07867_));
 OAI21_X1 _32850_ (.A(_05774_),
    .B1(_05834_),
    .B2(_05913_),
    .ZN(_07868_));
 NAND2_X1 _32851_ (.A1(_05774_),
    .A2(_07163_),
    .ZN(_07869_));
 NAND3_X1 _32852_ (.A1(_05807_),
    .A2(_05848_),
    .A3(_05749_),
    .ZN(_07870_));
 NAND4_X1 _32853_ (.A1(_07868_),
    .A2(_07869_),
    .A3(_07545_),
    .A4(_07870_),
    .ZN(_07871_));
 NAND2_X1 _32854_ (.A1(_06575_),
    .A2(_05751_),
    .ZN(_07873_));
 OAI21_X1 _32855_ (.A(_07873_),
    .B1(_05766_),
    .B2(_06646_),
    .ZN(_07874_));
 AND3_X1 _32856_ (.A1(_05751_),
    .A2(_05977_),
    .A3(_05763_),
    .ZN(_07875_));
 NOR4_X1 _32857_ (.A1(_07871_),
    .A2(_07187_),
    .A3(_07874_),
    .A4(_07875_),
    .ZN(_07876_));
 NAND3_X1 _32858_ (.A1(_05886_),
    .A2(_06662_),
    .A3(_05892_),
    .ZN(_07877_));
 OAI21_X1 _32859_ (.A(_06561_),
    .B1(_07156_),
    .B2(_05779_),
    .ZN(_07878_));
 OAI211_X1 _32860_ (.A(_06561_),
    .B(_05872_),
    .C1(_05851_),
    .C2(_05892_),
    .ZN(_07879_));
 OAI21_X1 _32861_ (.A(_05886_),
    .B1(_05834_),
    .B2(_06609_),
    .ZN(_07880_));
 AND4_X1 _32862_ (.A1(_07877_),
    .A2(_07878_),
    .A3(_07879_),
    .A4(_07880_),
    .ZN(_07881_));
 NAND4_X1 _32863_ (.A1(_07860_),
    .A2(_07867_),
    .A3(_07876_),
    .A4(_07881_),
    .ZN(_07882_));
 NOR2_X2 _32864_ (.A1(_07853_),
    .A2(_07882_),
    .ZN(_07884_));
 XOR2_X1 _32865_ (.A(_07884_),
    .B(_07478_),
    .Z(_07885_));
 XNOR2_X1 _32866_ (.A(_07827_),
    .B(_07885_),
    .ZN(_07886_));
 MUX2_X1 _32867_ (.A(_07632_),
    .B(_07886_),
    .S(_05069_),
    .Z(_00705_));
 XOR2_X1 _32868_ (.A(_17127_),
    .B(_16938_),
    .Z(_07887_));
 OAI21_X1 _32869_ (.A(_06384_),
    .B1(_05252_),
    .B2(_05301_),
    .ZN(_07888_));
 OAI21_X1 _32870_ (.A(_06384_),
    .B1(_05370_),
    .B2(_05332_),
    .ZN(_07889_));
 NAND3_X1 _32871_ (.A1(_07888_),
    .A2(_07889_),
    .A3(_07245_),
    .ZN(_07890_));
 NOR3_X1 _32872_ (.A1(_05384_),
    .A2(_05261_),
    .A3(_05389_),
    .ZN(_07891_));
 NOR2_X1 _32873_ (.A1(_07891_),
    .A2(_05381_),
    .ZN(_07892_));
 AOI211_X1 _32874_ (.A(_05164_),
    .B(_05274_),
    .C1(_07239_),
    .C2(_05257_),
    .ZN(_07894_));
 OAI211_X1 _32875_ (.A(_05353_),
    .B(_05172_),
    .C1(_05135_),
    .C2(_05150_),
    .ZN(_07895_));
 NAND2_X1 _32876_ (.A1(_05328_),
    .A2(_05142_),
    .ZN(_07896_));
 OAI211_X1 _32877_ (.A(_07895_),
    .B(_07896_),
    .C1(_05399_),
    .C2(_05432_),
    .ZN(_07897_));
 AOI21_X1 _32878_ (.A(_05274_),
    .B1(_07440_),
    .B2(_05433_),
    .ZN(_07898_));
 NOR4_X1 _32879_ (.A1(_07892_),
    .A2(_07894_),
    .A3(_07897_),
    .A4(_07898_),
    .ZN(_07899_));
 AOI22_X1 _32880_ (.A1(_05127_),
    .A2(_05353_),
    .B1(_05316_),
    .B2(_05143_),
    .ZN(_07900_));
 AND3_X1 _32881_ (.A1(_05413_),
    .A2(_06427_),
    .A3(_07900_),
    .ZN(_07901_));
 INV_X1 _32882_ (.A(_07266_),
    .ZN(_07902_));
 OAI211_X1 _32883_ (.A(_05180_),
    .B(_05206_),
    .C1(_06394_),
    .C2(_05438_),
    .ZN(_07903_));
 AND4_X1 _32884_ (.A1(_06403_),
    .A2(_06760_),
    .A3(_07902_),
    .A4(_07903_),
    .ZN(_07905_));
 AOI22_X1 _32885_ (.A1(_05248_),
    .A2(_05328_),
    .B1(_05209_),
    .B2(_05131_),
    .ZN(_07906_));
 AOI22_X1 _32886_ (.A1(_05260_),
    .A2(_05198_),
    .B1(_05243_),
    .B2(_05316_),
    .ZN(_07907_));
 AND4_X1 _32887_ (.A1(_05308_),
    .A2(_05305_),
    .A3(_07906_),
    .A4(_07907_),
    .ZN(_07908_));
 NAND4_X1 _32888_ (.A1(_07899_),
    .A2(_07901_),
    .A3(_07905_),
    .A4(_07908_),
    .ZN(_07909_));
 NAND2_X1 _32889_ (.A1(_07725_),
    .A2(_05281_),
    .ZN(_07910_));
 NAND3_X1 _32890_ (.A1(_05477_),
    .A2(_05449_),
    .A3(_05436_),
    .ZN(_07911_));
 OAI21_X1 _32891_ (.A(_05297_),
    .B1(_07911_),
    .B2(_05312_),
    .ZN(_07912_));
 NOR4_X1 _32892_ (.A1(_05193_),
    .A2(_05284_),
    .A3(_05312_),
    .A4(_05462_),
    .ZN(_07913_));
 OAI211_X1 _32893_ (.A(_07910_),
    .B(_07912_),
    .C1(_05342_),
    .C2(_07913_),
    .ZN(_07914_));
 AND2_X1 _32894_ (.A1(_05250_),
    .A2(_05353_),
    .ZN(_07916_));
 AOI22_X1 _32895_ (.A1(_05232_),
    .A2(_05347_),
    .B1(_05353_),
    .B2(_05141_),
    .ZN(_07917_));
 OAI221_X1 _32896_ (.A(_07917_),
    .B1(_05477_),
    .B2(_05255_),
    .C1(_05273_),
    .C2(_05432_),
    .ZN(_07918_));
 AND2_X1 _32897_ (.A1(_05198_),
    .A2(_05232_),
    .ZN(_07919_));
 OR2_X1 _32898_ (.A1(_07919_),
    .A2(_05471_),
    .ZN(_07920_));
 OR2_X1 _32899_ (.A1(_05422_),
    .A2(_05132_),
    .ZN(_07921_));
 OR4_X1 _32900_ (.A1(_07916_),
    .A2(_07918_),
    .A3(_07920_),
    .A4(_07921_),
    .ZN(_07922_));
 OR4_X1 _32901_ (.A1(_07890_),
    .A2(_07909_),
    .A3(_07914_),
    .A4(_07922_),
    .ZN(_07923_));
 OAI221_X1 _32902_ (.A(_05460_),
    .B1(_05294_),
    .B2(_05154_),
    .C1(_05273_),
    .C2(_05381_),
    .ZN(_07924_));
 AOI221_X4 _32903_ (.A(_07924_),
    .B1(_05248_),
    .B2(_06354_),
    .C1(_05389_),
    .C2(_05311_),
    .ZN(_07925_));
 AOI21_X1 _32904_ (.A(_06374_),
    .B1(_05295_),
    .B2(_05158_),
    .ZN(_07927_));
 AND3_X1 _32905_ (.A1(_05359_),
    .A2(_06394_),
    .A3(_05151_),
    .ZN(_07928_));
 NAND2_X1 _32906_ (.A1(_05199_),
    .A2(_05142_),
    .ZN(_07929_));
 OAI21_X1 _32907_ (.A(_07929_),
    .B1(_05339_),
    .B2(_07199_),
    .ZN(_07930_));
 NOR4_X1 _32908_ (.A1(_06805_),
    .A2(_07927_),
    .A3(_07928_),
    .A4(_07930_),
    .ZN(_07931_));
 AND2_X1 _32909_ (.A1(_05407_),
    .A2(_06354_),
    .ZN(_07932_));
 NOR4_X1 _32910_ (.A1(_07932_),
    .A2(_07738_),
    .A3(_06788_),
    .A4(_07265_),
    .ZN(_07933_));
 OAI21_X1 _32911_ (.A(_05220_),
    .B1(_07237_),
    .B2(_05237_),
    .ZN(_07934_));
 NAND3_X1 _32912_ (.A1(_05220_),
    .A2(_05348_),
    .A3(_05343_),
    .ZN(_07935_));
 NAND4_X1 _32913_ (.A1(_05215_),
    .A2(_06410_),
    .A3(_05172_),
    .A4(_05267_),
    .ZN(_07936_));
 AND4_X1 _32914_ (.A1(_05367_),
    .A2(_07934_),
    .A3(_07935_),
    .A4(_07936_),
    .ZN(_07938_));
 NAND4_X1 _32915_ (.A1(_07925_),
    .A2(_07931_),
    .A3(_07933_),
    .A4(_07938_),
    .ZN(_07939_));
 NOR2_X2 _32916_ (.A1(_07923_),
    .A2(_07939_),
    .ZN(_07940_));
 AND4_X1 _32917_ (.A1(_05567_),
    .A2(_05638_),
    .A3(_05535_),
    .A4(_05561_),
    .ZN(_07941_));
 AND2_X1 _32918_ (.A1(_05662_),
    .A2(_05584_),
    .ZN(_07942_));
 AOI211_X1 _32919_ (.A(_07941_),
    .B(_07942_),
    .C1(_07327_),
    .C2(_05670_),
    .ZN(_07943_));
 OAI21_X1 _32920_ (.A(_05670_),
    .B1(_05703_),
    .B2(_05705_),
    .ZN(_07944_));
 AND3_X1 _32921_ (.A1(_07943_),
    .A2(_07656_),
    .A3(_07944_),
    .ZN(_07945_));
 AOI211_X1 _32922_ (.A(_06263_),
    .B(_05652_),
    .C1(_05515_),
    .C2(_05593_),
    .ZN(_07946_));
 AND3_X1 _32923_ (.A1(_05651_),
    .A2(_05664_),
    .A3(_05686_),
    .ZN(_07947_));
 AND4_X1 _32924_ (.A1(_05593_),
    .A2(_06312_),
    .A3(_05525_),
    .A4(_05716_),
    .ZN(_07949_));
 AND4_X1 _32925_ (.A1(_05593_),
    .A2(_05638_),
    .A3(_06285_),
    .A4(_05716_),
    .ZN(_07950_));
 NOR4_X1 _32926_ (.A1(_07946_),
    .A2(_07947_),
    .A3(_07949_),
    .A4(_07950_),
    .ZN(_07951_));
 AOI21_X1 _32927_ (.A(_05649_),
    .B1(_06261_),
    .B2(_06704_),
    .ZN(_07952_));
 AOI211_X1 _32928_ (.A(_06298_),
    .B(_07952_),
    .C1(_05657_),
    .C2(_06299_),
    .ZN(_07953_));
 NAND2_X1 _32929_ (.A1(_05673_),
    .A2(_06346_),
    .ZN(_07954_));
 NOR2_X1 _32930_ (.A1(_05675_),
    .A2(_07285_),
    .ZN(_07955_));
 OR2_X1 _32931_ (.A1(_06319_),
    .A2(_05539_),
    .ZN(_07956_));
 NAND2_X1 _32932_ (.A1(_05672_),
    .A2(_06268_),
    .ZN(_07957_));
 AND4_X1 _32933_ (.A1(_07954_),
    .A2(_07955_),
    .A3(_07956_),
    .A4(_07957_),
    .ZN(_07958_));
 AND4_X1 _32934_ (.A1(_07945_),
    .A2(_07951_),
    .A3(_07953_),
    .A4(_07958_),
    .ZN(_07960_));
 OAI21_X1 _32935_ (.A(_05541_),
    .B1(_05690_),
    .B2(_05521_),
    .ZN(_07961_));
 OAI21_X1 _32936_ (.A(_05541_),
    .B1(_07301_),
    .B2(_06346_),
    .ZN(_07962_));
 AND3_X1 _32937_ (.A1(_07961_),
    .A2(_07962_),
    .A3(_07319_),
    .ZN(_07963_));
 AND3_X1 _32938_ (.A1(_05575_),
    .A2(_05506_),
    .A3(_05596_),
    .ZN(_07964_));
 NAND2_X1 _32939_ (.A1(_05547_),
    .A2(_05521_),
    .ZN(_07965_));
 NAND2_X1 _32940_ (.A1(_05646_),
    .A2(_05554_),
    .ZN(_07966_));
 NAND2_X1 _32941_ (.A1(_07965_),
    .A2(_07966_),
    .ZN(_07967_));
 AOI211_X1 _32942_ (.A(_07964_),
    .B(_07967_),
    .C1(_05703_),
    .C2(_05554_),
    .ZN(_07968_));
 INV_X1 _32943_ (.A(_07365_),
    .ZN(_07969_));
 NOR4_X1 _32944_ (.A1(_06752_),
    .A2(_07969_),
    .A3(_07633_),
    .A4(_05523_),
    .ZN(_07971_));
 AND2_X1 _32945_ (.A1(_05557_),
    .A2(_06251_),
    .ZN(_07972_));
 AND2_X1 _32946_ (.A1(_05562_),
    .A2(_05601_),
    .ZN(_07973_));
 NOR4_X1 _32947_ (.A1(_07683_),
    .A2(_05571_),
    .A3(_07972_),
    .A4(_07973_),
    .ZN(_07974_));
 AND4_X1 _32948_ (.A1(_07963_),
    .A2(_07968_),
    .A3(_07971_),
    .A4(_07974_),
    .ZN(_07975_));
 OAI21_X1 _32949_ (.A(_05583_),
    .B1(_05701_),
    .B2(_07324_),
    .ZN(_07976_));
 NAND3_X1 _32950_ (.A1(_05534_),
    .A2(_05583_),
    .A3(_05537_),
    .ZN(_07977_));
 AND2_X1 _32951_ (.A1(_07976_),
    .A2(_07977_),
    .ZN(_07978_));
 AOI21_X1 _32952_ (.A(_05598_),
    .B1(_06703_),
    .B2(_05585_),
    .ZN(_07979_));
 AND2_X1 _32953_ (.A1(_05606_),
    .A2(_05690_),
    .ZN(_07980_));
 AND4_X1 _32954_ (.A1(_05589_),
    .A2(_05596_),
    .A3(_06273_),
    .A4(_05572_),
    .ZN(_07982_));
 NOR4_X1 _32955_ (.A1(_07979_),
    .A2(_05600_),
    .A3(_07980_),
    .A4(_07982_),
    .ZN(_07983_));
 AND2_X1 _32956_ (.A1(_07330_),
    .A2(_05625_),
    .ZN(_07984_));
 AND2_X1 _32957_ (.A1(_06275_),
    .A2(_05626_),
    .ZN(_07985_));
 AND2_X1 _32958_ (.A1(_05626_),
    .A2(_06267_),
    .ZN(_07986_));
 AND4_X1 _32959_ (.A1(_05590_),
    .A2(_06273_),
    .A3(_05567_),
    .A4(_05561_),
    .ZN(_07987_));
 NOR4_X1 _32960_ (.A1(_07984_),
    .A2(_07985_),
    .A3(_07986_),
    .A4(_07987_),
    .ZN(_07988_));
 OAI21_X1 _32961_ (.A(_06266_),
    .B1(_05624_),
    .B2(_05686_),
    .ZN(_07989_));
 AND3_X1 _32962_ (.A1(_07989_),
    .A2(_06277_),
    .A3(_07335_),
    .ZN(_07990_));
 AND4_X1 _32963_ (.A1(_07978_),
    .A2(_07983_),
    .A3(_07988_),
    .A4(_07990_),
    .ZN(_07991_));
 OAI21_X1 _32964_ (.A(_05722_),
    .B1(_07668_),
    .B2(_05534_),
    .ZN(_07993_));
 OAI21_X1 _32965_ (.A(_06711_),
    .B1(_06267_),
    .B2(_05646_),
    .ZN(_07994_));
 NAND2_X1 _32966_ (.A1(_05710_),
    .A2(_05704_),
    .ZN(_07995_));
 NAND4_X1 _32967_ (.A1(_06285_),
    .A2(_05713_),
    .A3(_05714_),
    .A4(_05716_),
    .ZN(_07996_));
 AND4_X1 _32968_ (.A1(_06332_),
    .A2(_07994_),
    .A3(_07995_),
    .A4(_07996_),
    .ZN(_07997_));
 OAI21_X1 _32969_ (.A(_05696_),
    .B1(_05701_),
    .B2(_07324_),
    .ZN(_07998_));
 NAND4_X1 _32970_ (.A1(_05686_),
    .A2(_06272_),
    .A3(_05714_),
    .A4(_05666_),
    .ZN(_07999_));
 NAND4_X1 _32971_ (.A1(_06272_),
    .A2(_06291_),
    .A3(_05593_),
    .A4(_05714_),
    .ZN(_08000_));
 AND3_X1 _32972_ (.A1(_07998_),
    .A2(_07999_),
    .A3(_08000_),
    .ZN(_08001_));
 NAND2_X1 _32973_ (.A1(_05690_),
    .A2(_06343_),
    .ZN(_08002_));
 NAND2_X1 _32974_ (.A1(_05633_),
    .A2(_06343_),
    .ZN(_08004_));
 NAND2_X1 _32975_ (.A1(_06343_),
    .A2(_05616_),
    .ZN(_08005_));
 AND4_X1 _32976_ (.A1(_08002_),
    .A2(_06702_),
    .A3(_08004_),
    .A4(_08005_),
    .ZN(_08006_));
 AND4_X1 _32977_ (.A1(_07993_),
    .A2(_07997_),
    .A3(_08001_),
    .A4(_08006_),
    .ZN(_08007_));
 NAND4_X1 _32978_ (.A1(_07960_),
    .A2(_07975_),
    .A3(_07991_),
    .A4(_08007_),
    .ZN(_08008_));
 NOR2_X2 _32979_ (.A1(_08008_),
    .A2(_05733_),
    .ZN(_08009_));
 XOR2_X2 _32980_ (.A(_07940_),
    .B(_08009_),
    .Z(_08010_));
 AND4_X1 _32981_ (.A1(_06043_),
    .A2(_06213_),
    .A3(_06150_),
    .A4(_06183_),
    .ZN(_08011_));
 AND2_X1 _32982_ (.A1(_07081_),
    .A2(_06143_),
    .ZN(_08012_));
 AOI211_X1 _32983_ (.A(_08011_),
    .B(_08012_),
    .C1(_06041_),
    .C2(_07081_),
    .ZN(_08013_));
 OAI21_X1 _32984_ (.A(_07081_),
    .B1(_06107_),
    .B2(_06052_),
    .ZN(_08015_));
 OAI21_X1 _32985_ (.A(_07081_),
    .B1(_06099_),
    .B2(_06482_),
    .ZN(_08016_));
 AND3_X1 _32986_ (.A1(_08013_),
    .A2(_08015_),
    .A3(_08016_),
    .ZN(_08017_));
 AND2_X1 _32987_ (.A1(_06023_),
    .A2(_06170_),
    .ZN(_08018_));
 AND3_X1 _32988_ (.A1(_06190_),
    .A2(_06021_),
    .A3(_06213_),
    .ZN(_08019_));
 OR3_X1 _32989_ (.A1(_07761_),
    .A2(_08018_),
    .A3(_08019_),
    .ZN(_08020_));
 NAND2_X1 _32990_ (.A1(_06145_),
    .A2(_06869_),
    .ZN(_08021_));
 OAI21_X1 _32991_ (.A(_08021_),
    .B1(_06174_),
    .B2(_06176_),
    .ZN(_08022_));
 AND3_X1 _32992_ (.A1(_06180_),
    .A2(_06007_),
    .A3(_06150_),
    .ZN(_08023_));
 NOR4_X1 _32993_ (.A1(_08020_),
    .A2(_06840_),
    .A3(_08022_),
    .A4(_08023_),
    .ZN(_08024_));
 INV_X1 _32994_ (.A(_06517_),
    .ZN(_08026_));
 OR2_X1 _32995_ (.A1(_06120_),
    .A2(_06509_),
    .ZN(_08027_));
 AND4_X1 _32996_ (.A1(_06533_),
    .A2(_08026_),
    .A3(_08027_),
    .A4(_07074_),
    .ZN(_08028_));
 OAI21_X1 _32997_ (.A(_06224_),
    .B1(_07070_),
    .B2(_06484_),
    .ZN(_08029_));
 NAND3_X1 _32998_ (.A1(_06197_),
    .A2(_06125_),
    .A3(_06059_),
    .ZN(_08030_));
 AND3_X1 _32999_ (.A1(_07569_),
    .A2(_08029_),
    .A3(_08030_),
    .ZN(_08031_));
 AND2_X1 _33000_ (.A1(_06153_),
    .A2(_06052_),
    .ZN(_08032_));
 AND2_X1 _33001_ (.A1(_06844_),
    .A2(_06091_),
    .ZN(_08033_));
 NOR4_X1 _33002_ (.A1(_08032_),
    .A2(_08033_),
    .A3(_07063_),
    .A4(_07788_),
    .ZN(_08034_));
 AND4_X1 _33003_ (.A1(_08024_),
    .A2(_08028_),
    .A3(_08031_),
    .A4(_08034_),
    .ZN(_08035_));
 NAND3_X1 _33004_ (.A1(_07034_),
    .A2(_07030_),
    .A3(_06868_),
    .ZN(_08037_));
 AOI21_X1 _33005_ (.A(_06464_),
    .B1(_06458_),
    .B2(_07606_),
    .ZN(_08038_));
 AOI21_X1 _33006_ (.A(_06464_),
    .B1(_07782_),
    .B2(_07783_),
    .ZN(_08039_));
 NOR4_X1 _33007_ (.A1(_08037_),
    .A2(_06232_),
    .A3(_08038_),
    .A4(_08039_),
    .ZN(_08040_));
 NAND2_X1 _33008_ (.A1(_06038_),
    .A2(_06168_),
    .ZN(_08041_));
 NAND4_X1 _33009_ (.A1(_06892_),
    .A2(_06549_),
    .A3(_08041_),
    .A4(_06890_),
    .ZN(_08042_));
 OAI221_X1 _33010_ (.A(_06154_),
    .B1(_06467_),
    .B2(_06064_),
    .C1(_06042_),
    .C2(_06140_),
    .ZN(_08043_));
 NOR3_X1 _33011_ (.A1(_08042_),
    .A2(_08043_),
    .A3(_06129_),
    .ZN(_08044_));
 AND4_X1 _33012_ (.A1(_08017_),
    .A2(_08035_),
    .A3(_08040_),
    .A4(_08044_),
    .ZN(_08045_));
 AOI221_X4 _33013_ (.A(_07807_),
    .B1(_06086_),
    .B2(_06035_),
    .C1(_06041_),
    .C2(_06082_),
    .ZN(_08046_));
 OR4_X1 _33014_ (.A1(_06217_),
    .A2(_07041_),
    .A3(_07044_),
    .A4(_07024_),
    .ZN(_08048_));
 NAND2_X1 _33015_ (.A1(_06210_),
    .A2(_06049_),
    .ZN(_08049_));
 OAI21_X1 _33016_ (.A(_08049_),
    .B1(_06161_),
    .B2(_06851_),
    .ZN(_08050_));
 OAI22_X1 _33017_ (.A1(_06140_),
    .A2(_07783_),
    .B1(_06120_),
    .B2(_06851_),
    .ZN(_08051_));
 NOR4_X1 _33018_ (.A1(_08048_),
    .A2(_07101_),
    .A3(_08050_),
    .A4(_08051_),
    .ZN(_08052_));
 NAND3_X1 _33019_ (.A1(_06023_),
    .A2(_06484_),
    .A3(_06008_),
    .ZN(_08053_));
 NAND3_X1 _33020_ (.A1(_06889_),
    .A2(_07025_),
    .A3(_06065_),
    .ZN(_08054_));
 AND4_X1 _33021_ (.A1(_06909_),
    .A2(_08053_),
    .A3(_06870_),
    .A4(_08054_),
    .ZN(_08055_));
 NOR3_X1 _33022_ (.A1(_06164_),
    .A2(_06543_),
    .A3(_06462_),
    .ZN(_08056_));
 AOI22_X1 _33023_ (.A1(_06482_),
    .A2(_06849_),
    .B1(_06170_),
    .B2(_07025_),
    .ZN(_08057_));
 AOI22_X1 _33024_ (.A1(_06107_),
    .A2(_06137_),
    .B1(_06849_),
    .B2(_06076_),
    .ZN(_08059_));
 AND4_X1 _33025_ (.A1(_08055_),
    .A2(_08056_),
    .A3(_08057_),
    .A4(_08059_),
    .ZN(_08060_));
 OAI21_X1 _33026_ (.A(_06111_),
    .B1(_06076_),
    .B2(_06151_),
    .ZN(_08061_));
 OAI21_X1 _33027_ (.A(_08061_),
    .B1(_06458_),
    .B2(_06539_),
    .ZN(_08062_));
 NOR2_X1 _33028_ (.A1(_06866_),
    .A2(_06230_),
    .ZN(_08063_));
 AND2_X1 _33029_ (.A1(_06844_),
    .A2(_06223_),
    .ZN(_08064_));
 AOI21_X1 _33030_ (.A(_06088_),
    .B1(_07782_),
    .B2(_06872_),
    .ZN(_08065_));
 NOR4_X1 _33031_ (.A1(_08062_),
    .A2(_08063_),
    .A3(_08064_),
    .A4(_08065_),
    .ZN(_08066_));
 AND4_X1 _33032_ (.A1(_08046_),
    .A2(_08052_),
    .A3(_08060_),
    .A4(_08066_),
    .ZN(_08067_));
 NAND2_X2 _33033_ (.A1(_08045_),
    .A2(_08067_),
    .ZN(_08068_));
 XNOR2_X1 _33034_ (.A(_08068_),
    .B(_00995_),
    .ZN(_08070_));
 XNOR2_X1 _33035_ (.A(_08010_),
    .B(_08070_),
    .ZN(_08071_));
 OR4_X1 _33036_ (.A1(_06593_),
    .A2(_06976_),
    .A3(_07003_),
    .A4(_06995_),
    .ZN(_08072_));
 OAI211_X1 _33037_ (.A(_05971_),
    .B(_07873_),
    .C1(_06646_),
    .C2(_07155_),
    .ZN(_08073_));
 AOI22_X1 _33038_ (.A1(_05857_),
    .A2(_05974_),
    .B1(_05958_),
    .B2(_07163_),
    .ZN(_08074_));
 OAI221_X1 _33039_ (.A(_08074_),
    .B1(_07500_),
    .B2(_07113_),
    .C1(_06591_),
    .C2(_06569_),
    .ZN(_08075_));
 NOR4_X1 _33040_ (.A1(_08072_),
    .A2(_06654_),
    .A3(_08073_),
    .A4(_08075_),
    .ZN(_08076_));
 INV_X1 _33041_ (.A(_06608_),
    .ZN(_08077_));
 INV_X1 _33042_ (.A(_07528_),
    .ZN(_08078_));
 AOI21_X1 _33043_ (.A(_06960_),
    .B1(_08077_),
    .B2(_08078_),
    .ZN(_08079_));
 INV_X1 _33044_ (.A(_05861_),
    .ZN(_08081_));
 AOI21_X1 _33045_ (.A(_08081_),
    .B1(_06961_),
    .B2(_06997_),
    .ZN(_08082_));
 AND3_X1 _33046_ (.A1(_05974_),
    .A2(_05872_),
    .A3(_05851_),
    .ZN(_08083_));
 NOR4_X1 _33047_ (.A1(_08079_),
    .A2(_08082_),
    .A3(_07168_),
    .A4(_08083_),
    .ZN(_08084_));
 NAND2_X1 _33048_ (.A1(_05952_),
    .A2(_05937_),
    .ZN(_08085_));
 NAND2_X1 _33049_ (.A1(_05856_),
    .A2(_05827_),
    .ZN(_08086_));
 NAND2_X1 _33050_ (.A1(_08085_),
    .A2(_08086_),
    .ZN(_08087_));
 AOI221_X4 _33051_ (.A(_08087_),
    .B1(_05763_),
    .B2(_07005_),
    .C1(_05807_),
    .C2(_05909_),
    .ZN(_08088_));
 OAI21_X1 _33052_ (.A(_07010_),
    .B1(_05766_),
    .B2(_06598_),
    .ZN(_08089_));
 AOI221_X4 _33053_ (.A(_08089_),
    .B1(_05967_),
    .B2(_05807_),
    .C1(_05771_),
    .C2(_05959_),
    .ZN(_08090_));
 OAI21_X1 _33054_ (.A(_05912_),
    .B1(_05817_),
    .B2(_05864_),
    .ZN(_08092_));
 AOI22_X1 _33055_ (.A1(_05974_),
    .A2(_05817_),
    .B1(_05773_),
    .B2(_05886_),
    .ZN(_08093_));
 AND4_X1 _33056_ (.A1(_08088_),
    .A2(_08090_),
    .A3(_08092_),
    .A4(_08093_),
    .ZN(_08094_));
 AOI21_X1 _33057_ (.A(_06643_),
    .B1(_06607_),
    .B2(_07155_),
    .ZN(_08095_));
 NOR2_X1 _33058_ (.A1(_08095_),
    .A2(_07549_),
    .ZN(_08096_));
 OAI21_X1 _33059_ (.A(_05958_),
    .B1(_05955_),
    .B2(_05844_),
    .ZN(_08097_));
 OAI21_X1 _33060_ (.A(_06561_),
    .B1(_05913_),
    .B2(_05977_),
    .ZN(_08098_));
 AND4_X1 _33061_ (.A1(_07016_),
    .A2(_08096_),
    .A3(_08097_),
    .A4(_08098_),
    .ZN(_08099_));
 AND4_X1 _33062_ (.A1(_08076_),
    .A2(_08084_),
    .A3(_08094_),
    .A4(_08099_),
    .ZN(_08100_));
 OAI21_X1 _33063_ (.A(_05793_),
    .B1(_06566_),
    .B2(_06569_),
    .ZN(_08101_));
 AOI21_X1 _33064_ (.A(_08101_),
    .B1(_05774_),
    .B2(_06605_),
    .ZN(_08103_));
 AOI21_X1 _33065_ (.A(_06598_),
    .B1(_07500_),
    .B2(_06970_),
    .ZN(_08104_));
 AND2_X1 _33066_ (.A1(_05972_),
    .A2(_06609_),
    .ZN(_08105_));
 AND2_X1 _33067_ (.A1(_05979_),
    .A2(_05794_),
    .ZN(_08106_));
 NOR3_X1 _33068_ (.A1(_08104_),
    .A2(_08105_),
    .A3(_08106_),
    .ZN(_08107_));
 AND4_X1 _33069_ (.A1(_06658_),
    .A2(_08103_),
    .A3(_06659_),
    .A4(_08107_),
    .ZN(_08108_));
 AND2_X1 _33070_ (.A1(_05864_),
    .A2(_05803_),
    .ZN(_08109_));
 OR4_X1 _33071_ (.A1(_05943_),
    .A2(_05926_),
    .A3(_05932_),
    .A4(_08109_),
    .ZN(_08110_));
 NAND3_X1 _33072_ (.A1(_05751_),
    .A2(_06572_),
    .A3(_05779_),
    .ZN(_08111_));
 OAI211_X1 _33073_ (.A(_05914_),
    .B(_08111_),
    .C1(_05812_),
    .C2(_05922_),
    .ZN(_08112_));
 OR2_X1 _33074_ (.A1(_05815_),
    .A2(_05904_),
    .ZN(_08114_));
 NOR4_X1 _33075_ (.A1(_08110_),
    .A2(_05772_),
    .A3(_08112_),
    .A4(_08114_),
    .ZN(_08115_));
 NOR4_X1 _33076_ (.A1(_06942_),
    .A2(_06631_),
    .A3(_06634_),
    .A4(_07152_),
    .ZN(_08116_));
 NAND2_X1 _33077_ (.A1(_05876_),
    .A2(_05809_),
    .ZN(_08117_));
 AOI22_X1 _33078_ (.A1(_06604_),
    .A2(_05831_),
    .B1(_05828_),
    .B2(_06595_),
    .ZN(_08118_));
 AND4_X1 _33079_ (.A1(_07496_),
    .A2(_08116_),
    .A3(_08117_),
    .A4(_08118_),
    .ZN(_08119_));
 AND2_X1 _33080_ (.A1(_06609_),
    .A2(_05886_),
    .ZN(_08120_));
 AND3_X1 _33081_ (.A1(_05867_),
    .A2(_05849_),
    .A3(_05825_),
    .ZN(_08121_));
 NOR4_X1 _33082_ (.A1(_07524_),
    .A2(_07830_),
    .A3(_08120_),
    .A4(_08121_),
    .ZN(_08122_));
 AND4_X1 _33083_ (.A1(_08108_),
    .A2(_08115_),
    .A3(_08119_),
    .A4(_08122_),
    .ZN(_08123_));
 NAND2_X2 _33084_ (.A1(_08100_),
    .A2(_08123_),
    .ZN(_08125_));
 XNOR2_X1 _33085_ (.A(_08125_),
    .B(_07756_),
    .ZN(_08126_));
 XNOR2_X1 _33086_ (.A(_08071_),
    .B(_08126_),
    .ZN(_08127_));
 MUX2_X1 _33087_ (.A(_07887_),
    .B(_08127_),
    .S(_05069_),
    .Z(_00706_));
 XOR2_X1 _33088_ (.A(_17128_),
    .B(_16939_),
    .Z(_08128_));
 AOI211_X1 _33089_ (.A(_05685_),
    .B(_05682_),
    .C1(_05515_),
    .C2(_16719_),
    .ZN(_08129_));
 AND2_X1 _33090_ (.A1(_05534_),
    .A2(_05681_),
    .ZN(_08130_));
 OR4_X1 _33091_ (.A1(_05684_),
    .A2(_08129_),
    .A3(_06339_),
    .A4(_08130_),
    .ZN(_08131_));
 AND2_X1 _33092_ (.A1(_05721_),
    .A2(_07339_),
    .ZN(_08132_));
 AOI21_X1 _33093_ (.A(_07649_),
    .B1(_06675_),
    .B2(_05549_),
    .ZN(_08133_));
 NOR4_X1 _33094_ (.A1(_08131_),
    .A2(_07302_),
    .A3(_08132_),
    .A4(_08133_),
    .ZN(_08135_));
 NAND3_X1 _33095_ (.A1(_05644_),
    .A2(_06242_),
    .A3(_05679_),
    .ZN(_08136_));
 NAND2_X1 _33096_ (.A1(_08136_),
    .A2(_07404_),
    .ZN(_08137_));
 AND3_X1 _33097_ (.A1(_06271_),
    .A2(_05529_),
    .A3(_05679_),
    .ZN(_08138_));
 NOR3_X1 _33098_ (.A1(_08137_),
    .A2(_07295_),
    .A3(_08138_),
    .ZN(_08139_));
 OAI21_X1 _33099_ (.A(_05710_),
    .B1(_05534_),
    .B2(_06268_),
    .ZN(_08140_));
 OAI211_X1 _33100_ (.A(_05710_),
    .B(_05493_),
    .C1(_05515_),
    .C2(_05611_),
    .ZN(_08141_));
 AND4_X1 _33101_ (.A1(_07995_),
    .A2(_08139_),
    .A3(_08140_),
    .A4(_08141_),
    .ZN(_08142_));
 AND3_X1 _33102_ (.A1(_05704_),
    .A2(_05488_),
    .A3(_05637_),
    .ZN(_08143_));
 AND4_X1 _33103_ (.A1(_05524_),
    .A2(_05637_),
    .A3(_05498_),
    .A4(_05487_),
    .ZN(_08144_));
 OR3_X1 _33104_ (.A1(_07947_),
    .A2(_08143_),
    .A3(_08144_),
    .ZN(_08146_));
 AOI21_X1 _33105_ (.A(_05649_),
    .B1(_05602_),
    .B2(_06713_),
    .ZN(_08147_));
 AND3_X1 _33106_ (.A1(_05642_),
    .A2(_05664_),
    .A3(_06271_),
    .ZN(_08148_));
 NOR4_X1 _33107_ (.A1(_08146_),
    .A2(_07275_),
    .A3(_08147_),
    .A4(_08148_),
    .ZN(_08149_));
 NAND2_X1 _33108_ (.A1(_05672_),
    .A2(_05704_),
    .ZN(_08150_));
 OAI21_X1 _33109_ (.A(_05672_),
    .B1(_05605_),
    .B2(_05575_),
    .ZN(_08151_));
 NAND4_X1 _33110_ (.A1(_06690_),
    .A2(_08150_),
    .A3(_07957_),
    .A4(_08151_),
    .ZN(_08152_));
 NOR4_X1 _33111_ (.A1(_08152_),
    .A2(_07679_),
    .A3(_05669_),
    .A4(_07942_),
    .ZN(_08153_));
 AND4_X1 _33112_ (.A1(_08135_),
    .A2(_08142_),
    .A3(_08149_),
    .A4(_08153_),
    .ZN(_08154_));
 OAI21_X1 _33113_ (.A(_05609_),
    .B1(_06697_),
    .B2(_05570_),
    .ZN(_08155_));
 NAND4_X1 _33114_ (.A1(_06242_),
    .A2(_05581_),
    .A3(_16719_),
    .A4(_05514_),
    .ZN(_08157_));
 OAI21_X1 _33115_ (.A(_05608_),
    .B1(_05699_),
    .B2(_05564_),
    .ZN(_08158_));
 AND3_X1 _33116_ (.A1(_08155_),
    .A2(_08157_),
    .A3(_08158_),
    .ZN(_08159_));
 OAI21_X1 _33117_ (.A(_05582_),
    .B1(_06267_),
    .B2(_05645_),
    .ZN(_08160_));
 OAI21_X1 _33118_ (.A(_05582_),
    .B1(_05508_),
    .B2(_05692_),
    .ZN(_08161_));
 AND3_X1 _33119_ (.A1(_08159_),
    .A2(_08160_),
    .A3(_08161_),
    .ZN(_08162_));
 NAND4_X1 _33120_ (.A1(_06242_),
    .A2(_05496_),
    .A3(_05567_),
    .A4(_05486_),
    .ZN(_08163_));
 OAI211_X1 _33121_ (.A(_07655_),
    .B(_08163_),
    .C1(_06245_),
    .C2(_05585_),
    .ZN(_08164_));
 AOI211_X1 _33122_ (.A(_06263_),
    .B(_06245_),
    .C1(_05515_),
    .C2(_05590_),
    .ZN(_08165_));
 OAI211_X1 _33123_ (.A(_05490_),
    .B(_05493_),
    .C1(_05494_),
    .C2(_05590_),
    .ZN(_08166_));
 NAND4_X1 _33124_ (.A1(_05490_),
    .A2(_05657_),
    .A3(_05664_),
    .A4(_05524_),
    .ZN(_08168_));
 NAND2_X1 _33125_ (.A1(_08166_),
    .A2(_08168_),
    .ZN(_08169_));
 OAI21_X1 _33126_ (.A(_06243_),
    .B1(_06245_),
    .B2(_06249_),
    .ZN(_08170_));
 NOR4_X1 _33127_ (.A1(_08164_),
    .A2(_08165_),
    .A3(_08169_),
    .A4(_08170_),
    .ZN(_08171_));
 OAI21_X1 _33128_ (.A(_05597_),
    .B1(_07301_),
    .B2(_05558_),
    .ZN(_08172_));
 OAI21_X1 _33129_ (.A(_05597_),
    .B1(_05516_),
    .B2(_05616_),
    .ZN(_08173_));
 NAND3_X1 _33130_ (.A1(_08172_),
    .A2(_08173_),
    .A3(_06724_),
    .ZN(_08174_));
 AOI21_X1 _33131_ (.A(_06287_),
    .B1(_05658_),
    .B2(_05602_),
    .ZN(_08175_));
 NOR4_X1 _33132_ (.A1(_08174_),
    .A2(_08175_),
    .A3(_07984_),
    .A4(_07377_),
    .ZN(_08176_));
 NAND4_X1 _33133_ (.A1(_05551_),
    .A2(_05553_),
    .A3(_07965_),
    .A4(_07345_),
    .ZN(_08177_));
 AND2_X1 _33134_ (.A1(_05624_),
    .A2(_05562_),
    .ZN(_08179_));
 AOI21_X1 _33135_ (.A(_05563_),
    .B1(_05509_),
    .B2(_07650_),
    .ZN(_08180_));
 NOR4_X1 _33136_ (.A1(_08177_),
    .A2(_08179_),
    .A3(_07973_),
    .A4(_08180_),
    .ZN(_08181_));
 AND4_X1 _33137_ (.A1(_08162_),
    .A2(_08171_),
    .A3(_08176_),
    .A4(_08181_),
    .ZN(_08182_));
 AND2_X1 _33138_ (.A1(_08154_),
    .A2(_08182_),
    .ZN(_08183_));
 BUF_X2 _33139_ (.A(_08183_),
    .Z(_08184_));
 XNOR2_X2 _33140_ (.A(_08184_),
    .B(_05484_),
    .ZN(_08185_));
 AND2_X1 _33141_ (.A1(_06101_),
    .A2(_06119_),
    .ZN(_08186_));
 AND2_X1 _33142_ (.A1(_06102_),
    .A2(_06119_),
    .ZN(_08187_));
 AND2_X1 _33143_ (.A1(_06119_),
    .A2(_06143_),
    .ZN(_08188_));
 OR4_X1 _33144_ (.A1(_08186_),
    .A2(_06445_),
    .A3(_08187_),
    .A4(_08188_),
    .ZN(_08190_));
 OAI21_X1 _33145_ (.A(_06078_),
    .B1(_06869_),
    .B2(_07090_),
    .ZN(_08191_));
 OAI211_X1 _33146_ (.A(_06450_),
    .B(_08191_),
    .C1(_06088_),
    .C2(_06046_),
    .ZN(_08192_));
 NOR4_X1 _33147_ (.A1(_08190_),
    .A2(_08192_),
    .A3(_06121_),
    .A4(_06442_),
    .ZN(_08193_));
 AND3_X1 _33148_ (.A1(_06209_),
    .A2(_05992_),
    .A3(_06058_),
    .ZN(_08194_));
 OR4_X1 _33149_ (.A1(_06531_),
    .A2(_08194_),
    .A3(_07052_),
    .A4(_07761_),
    .ZN(_08195_));
 AND2_X1 _33150_ (.A1(_06482_),
    .A2(_07081_),
    .ZN(_08196_));
 AOI21_X1 _33151_ (.A(_06206_),
    .B1(_06851_),
    .B2(_06205_),
    .ZN(_08197_));
 NOR4_X1 _33152_ (.A1(_08195_),
    .A2(_07765_),
    .A3(_08196_),
    .A4(_08197_),
    .ZN(_08198_));
 AND2_X1 _33153_ (.A1(_06106_),
    .A2(_06110_),
    .ZN(_08199_));
 OR3_X1 _33154_ (.A1(_07024_),
    .A2(_08199_),
    .A3(_06453_),
    .ZN(_08201_));
 NAND2_X1 _33155_ (.A1(_06090_),
    .A2(_06211_),
    .ZN(_08202_));
 NAND3_X1 _33156_ (.A1(_07776_),
    .A2(_06471_),
    .A3(_08202_),
    .ZN(_08203_));
 AND2_X1 _33157_ (.A1(_06904_),
    .A2(_06045_),
    .ZN(_08204_));
 AOI21_X1 _33158_ (.A(_06117_),
    .B1(_06465_),
    .B2(_06455_),
    .ZN(_08205_));
 NOR4_X1 _33159_ (.A1(_08201_),
    .A2(_08203_),
    .A3(_08204_),
    .A4(_08205_),
    .ZN(_08206_));
 NAND2_X1 _33160_ (.A1(_06099_),
    .A2(_06221_),
    .ZN(_08207_));
 OAI21_X1 _33161_ (.A(_06197_),
    .B1(_06510_),
    .B2(_06522_),
    .ZN(_08208_));
 OAI21_X1 _33162_ (.A(_06197_),
    .B1(_06168_),
    .B2(_06466_),
    .ZN(_08209_));
 OAI21_X1 _33163_ (.A(_06221_),
    .B1(_06456_),
    .B2(_06101_),
    .ZN(_08210_));
 AND4_X1 _33164_ (.A1(_08207_),
    .A2(_08208_),
    .A3(_08209_),
    .A4(_08210_),
    .ZN(_08212_));
 AND4_X1 _33165_ (.A1(_08193_),
    .A2(_08198_),
    .A3(_08206_),
    .A4(_08212_),
    .ZN(_08213_));
 OAI211_X1 _33166_ (.A(_06063_),
    .B(_06058_),
    .C1(_06032_),
    .C2(_05986_),
    .ZN(_08214_));
 OAI21_X1 _33167_ (.A(_08214_),
    .B1(_06514_),
    .B2(_06064_),
    .ZN(_08215_));
 AOI21_X1 _33168_ (.A(_06040_),
    .B1(_07782_),
    .B2(_06054_),
    .ZN(_08216_));
 OAI21_X1 _33169_ (.A(_08041_),
    .B1(_06040_),
    .B2(_06046_),
    .ZN(_08217_));
 AOI21_X1 _33170_ (.A(_06064_),
    .B1(_06459_),
    .B2(_06467_),
    .ZN(_08218_));
 NOR4_X1 _33171_ (.A1(_08215_),
    .A2(_08216_),
    .A3(_08217_),
    .A4(_08218_),
    .ZN(_08219_));
 AOI211_X1 _33172_ (.A(_06491_),
    .B(_07103_),
    .C1(_07026_),
    .C2(_05997_),
    .ZN(_08220_));
 AND3_X1 _33173_ (.A1(_06103_),
    .A2(_06172_),
    .A3(_05993_),
    .ZN(_08221_));
 AOI211_X1 _33174_ (.A(_08221_),
    .B(_06486_),
    .C1(_06035_),
    .C2(_07026_),
    .ZN(_08223_));
 NOR4_X1 _33175_ (.A1(_06873_),
    .A2(_06483_),
    .A3(_06876_),
    .A4(_08018_),
    .ZN(_08224_));
 NAND4_X1 _33176_ (.A1(_08219_),
    .A2(_08220_),
    .A3(_08223_),
    .A4(_08224_),
    .ZN(_08225_));
 OAI21_X1 _33177_ (.A(_06844_),
    .B1(_05990_),
    .B2(_06521_),
    .ZN(_08226_));
 OAI21_X1 _33178_ (.A(_06844_),
    .B1(_06128_),
    .B2(_06151_),
    .ZN(_08227_));
 NAND3_X1 _33179_ (.A1(_08226_),
    .A2(_08227_),
    .A3(_06518_),
    .ZN(_08228_));
 AND3_X1 _33180_ (.A1(_06146_),
    .A2(_06021_),
    .A3(_06158_),
    .ZN(_08229_));
 AOI221_X4 _33181_ (.A(_08229_),
    .B1(_06466_),
    .B2(_06166_),
    .C1(_06044_),
    .C2(_07041_),
    .ZN(_08230_));
 NAND4_X1 _33182_ (.A1(_06521_),
    .A2(_06172_),
    .A3(_05987_),
    .A4(_06158_),
    .ZN(_08231_));
 OAI21_X1 _33183_ (.A(_06136_),
    .B1(_06075_),
    .B2(_06151_),
    .ZN(_08232_));
 OAI21_X1 _33184_ (.A(_06136_),
    .B1(_06482_),
    .B2(_06130_),
    .ZN(_08234_));
 AND2_X1 _33185_ (.A1(_08232_),
    .A2(_08234_),
    .ZN(_08235_));
 NAND4_X1 _33186_ (.A1(_08230_),
    .A2(_06173_),
    .A3(_08231_),
    .A4(_08235_),
    .ZN(_08236_));
 OAI211_X1 _33187_ (.A(_06037_),
    .B(_06158_),
    .C1(_06000_),
    .C2(_06143_),
    .ZN(_08237_));
 NAND4_X1 _33188_ (.A1(_08021_),
    .A2(_08237_),
    .A3(_07097_),
    .A4(_06152_),
    .ZN(_08238_));
 NOR4_X1 _33189_ (.A1(_08225_),
    .A2(_08228_),
    .A3(_08236_),
    .A4(_08238_),
    .ZN(_08239_));
 AND2_X1 _33190_ (.A1(_08213_),
    .A2(_08239_),
    .ZN(_08240_));
 BUF_X2 _33191_ (.A(_08240_),
    .Z(_08241_));
 XNOR2_X1 _33192_ (.A(_08241_),
    .B(_00996_),
    .ZN(_08242_));
 XNOR2_X1 _33193_ (.A(_08185_),
    .B(_08242_),
    .ZN(_08243_));
 OR4_X1 _33194_ (.A1(_05975_),
    .A2(_07485_),
    .A3(_08105_),
    .A4(_06937_),
    .ZN(_08245_));
 OAI21_X1 _33195_ (.A(_05958_),
    .B1(_05963_),
    .B2(_06977_),
    .ZN(_08246_));
 OAI211_X1 _33196_ (.A(_05948_),
    .B(_05748_),
    .C1(_05783_),
    .C2(_05794_),
    .ZN(_08247_));
 OAI211_X1 _33197_ (.A(_08246_),
    .B(_08247_),
    .C1(_06640_),
    .C2(_08078_),
    .ZN(_08248_));
 NAND4_X1 _33198_ (.A1(_07841_),
    .A2(_07133_),
    .A3(_07134_),
    .A4(_08085_),
    .ZN(_08249_));
 OAI211_X1 _33199_ (.A(_05979_),
    .B(_16802_),
    .C1(_05781_),
    .C2(_05737_),
    .ZN(_08250_));
 OAI211_X1 _33200_ (.A(_05948_),
    .B(_05802_),
    .C1(_07163_),
    .C2(_05829_),
    .ZN(_08251_));
 OAI211_X1 _33201_ (.A(_08250_),
    .B(_08251_),
    .C1(_08077_),
    .C2(_06591_),
    .ZN(_08252_));
 NOR4_X1 _33202_ (.A1(_08245_),
    .A2(_08248_),
    .A3(_08249_),
    .A4(_08252_),
    .ZN(_08253_));
 OAI21_X1 _33203_ (.A(_05751_),
    .B1(_06575_),
    .B2(_05892_),
    .ZN(_08254_));
 NAND2_X1 _33204_ (.A1(_06561_),
    .A2(_05866_),
    .ZN(_08256_));
 OAI211_X1 _33205_ (.A(_07558_),
    .B(_08256_),
    .C1(_05954_),
    .C2(_05871_),
    .ZN(_08257_));
 AND2_X1 _33206_ (.A1(_05870_),
    .A2(_05864_),
    .ZN(_08258_));
 OR2_X1 _33207_ (.A1(_08258_),
    .A2(_05877_),
    .ZN(_08259_));
 OAI211_X1 _33208_ (.A(_07010_),
    .B(_07560_),
    .C1(_05953_),
    .C2(_05890_),
    .ZN(_08260_));
 NOR4_X1 _33209_ (.A1(_08257_),
    .A2(_08259_),
    .A3(_05884_),
    .A4(_08260_),
    .ZN(_08261_));
 NAND2_X1 _33210_ (.A1(_05771_),
    .A2(_05834_),
    .ZN(_08262_));
 AND3_X1 _33211_ (.A1(_08262_),
    .A2(_07000_),
    .A3(_05784_),
    .ZN(_08263_));
 OAI21_X1 _33212_ (.A(_05774_),
    .B1(_05857_),
    .B2(_05807_),
    .ZN(_08264_));
 AND4_X1 _33213_ (.A1(_07544_),
    .A2(_08263_),
    .A3(_07545_),
    .A4(_08264_),
    .ZN(_08265_));
 AND4_X1 _33214_ (.A1(_08254_),
    .A2(_08261_),
    .A3(_07189_),
    .A4(_08265_),
    .ZN(_08267_));
 AND3_X1 _33215_ (.A1(_07550_),
    .A2(_07548_),
    .A3(_07856_),
    .ZN(_08268_));
 OAI211_X1 _33216_ (.A(_08268_),
    .B(_07551_),
    .C1(_06643_),
    .C2(_06987_),
    .ZN(_08269_));
 OAI21_X1 _33217_ (.A(_05861_),
    .B1(_05878_),
    .B2(_07528_),
    .ZN(_08270_));
 OAI21_X1 _33218_ (.A(_08270_),
    .B1(_08077_),
    .B2(_08081_),
    .ZN(_08271_));
 OAI21_X1 _33219_ (.A(_05828_),
    .B1(_07163_),
    .B2(_05829_),
    .ZN(_08272_));
 NAND2_X1 _33220_ (.A1(_05828_),
    .A2(_05811_),
    .ZN(_08273_));
 NAND2_X1 _33221_ (.A1(_05828_),
    .A2(_06559_),
    .ZN(_08274_));
 NAND4_X1 _33222_ (.A1(_08272_),
    .A2(_06661_),
    .A3(_08273_),
    .A4(_08274_),
    .ZN(_08275_));
 NAND2_X1 _33223_ (.A1(_05810_),
    .A2(_06571_),
    .ZN(_08276_));
 OR3_X1 _33224_ (.A1(_08276_),
    .A2(_05824_),
    .A3(_05818_),
    .ZN(_08278_));
 NOR4_X1 _33225_ (.A1(_08269_),
    .A2(_08271_),
    .A3(_08275_),
    .A4(_08278_),
    .ZN(_08279_));
 OAI21_X1 _33226_ (.A(_06604_),
    .B1(_05878_),
    .B2(_07528_),
    .ZN(_08280_));
 OAI211_X1 _33227_ (.A(_05848_),
    .B(_05906_),
    .C1(_07163_),
    .C2(_05937_),
    .ZN(_08281_));
 NAND4_X1 _33228_ (.A1(_05848_),
    .A2(_05892_),
    .A3(_05780_),
    .A4(_05906_),
    .ZN(_08282_));
 AND3_X1 _33229_ (.A1(_08280_),
    .A2(_08281_),
    .A3(_08282_),
    .ZN(_08283_));
 AND2_X1 _33230_ (.A1(_05931_),
    .A2(_05900_),
    .ZN(_08284_));
 NOR4_X1 _33231_ (.A1(_07123_),
    .A2(_05904_),
    .A3(_06628_),
    .A4(_08284_),
    .ZN(_08285_));
 INV_X1 _33232_ (.A(_05942_),
    .ZN(_08286_));
 NAND2_X1 _33233_ (.A1(_06559_),
    .A2(_05939_),
    .ZN(_08287_));
 OAI21_X1 _33234_ (.A(_05939_),
    .B1(_05807_),
    .B2(_05864_),
    .ZN(_08289_));
 AND4_X1 _33235_ (.A1(_08286_),
    .A2(_08287_),
    .A3(_07149_),
    .A4(_08289_),
    .ZN(_08290_));
 AOI21_X1 _33236_ (.A(_05922_),
    .B1(_07165_),
    .B2(_06569_),
    .ZN(_08291_));
 AOI21_X1 _33237_ (.A(_05922_),
    .B1(_06948_),
    .B2(_05769_),
    .ZN(_08292_));
 AOI211_X1 _33238_ (.A(_08291_),
    .B(_08292_),
    .C1(_05855_),
    .C2(_05912_),
    .ZN(_08293_));
 AND4_X1 _33239_ (.A1(_08283_),
    .A2(_08285_),
    .A3(_08290_),
    .A4(_08293_),
    .ZN(_08294_));
 NAND4_X1 _33240_ (.A1(_08253_),
    .A2(_08267_),
    .A3(_08279_),
    .A4(_08294_),
    .ZN(_08295_));
 NOR2_X2 _33241_ (.A1(_08295_),
    .A2(_07015_),
    .ZN(_08296_));
 XOR2_X1 _33242_ (.A(_07940_),
    .B(_08296_),
    .Z(_08297_));
 XNOR2_X1 _33243_ (.A(_08243_),
    .B(_08297_),
    .ZN(_08298_));
 BUF_X2 _33244_ (.A(_09038_),
    .Z(_08300_));
 MUX2_X1 _33245_ (.A(_08128_),
    .B(_08298_),
    .S(_08300_),
    .Z(_00707_));
 XOR2_X1 _33246_ (.A(_17129_),
    .B(_16940_),
    .Z(_08301_));
 XOR2_X1 _33247_ (.A(_06669_),
    .B(_00997_),
    .Z(_08302_));
 XOR2_X1 _33248_ (.A(_05734_),
    .B(_08241_),
    .Z(_08303_));
 XNOR2_X1 _33249_ (.A(_08303_),
    .B(_05369_),
    .ZN(_08304_));
 XNOR2_X1 _33250_ (.A(_08302_),
    .B(_08304_),
    .ZN(_08305_));
 MUX2_X1 _33251_ (.A(_08301_),
    .B(_08305_),
    .S(_08300_),
    .Z(_00668_));
 XOR2_X1 _33252_ (.A(_17130_),
    .B(_16941_),
    .Z(_08306_));
 INV_X1 _33253_ (.A(_08241_),
    .ZN(_08307_));
 XNOR2_X2 _33254_ (.A(_08307_),
    .B(_06233_),
    .ZN(_08309_));
 XNOR2_X1 _33255_ (.A(_06438_),
    .B(_08309_),
    .ZN(_08310_));
 XNOR2_X1 _33256_ (.A(_07017_),
    .B(_14977_),
    .ZN(_08311_));
 XNOR2_X1 _33257_ (.A(_08311_),
    .B(_06669_),
    .ZN(_08312_));
 XNOR2_X1 _33258_ (.A(_08310_),
    .B(_08312_),
    .ZN(_08313_));
 MUX2_X1 _33259_ (.A(_08306_),
    .B(_08313_),
    .S(_08300_),
    .Z(_00669_));
 XOR2_X1 _33260_ (.A(_17100_),
    .B(_16942_),
    .Z(_08314_));
 XOR2_X2 _33261_ (.A(_07017_),
    .B(_06553_),
    .Z(_08315_));
 XNOR2_X1 _33262_ (.A(_08315_),
    .B(_06836_),
    .ZN(_08316_));
 XNOR2_X1 _33263_ (.A(_07193_),
    .B(_00999_),
    .ZN(_08317_));
 XNOR2_X1 _33264_ (.A(_08316_),
    .B(_08317_),
    .ZN(_08319_));
 MUX2_X1 _33265_ (.A(_08314_),
    .B(_08319_),
    .S(_08300_),
    .Z(_00670_));
 XOR2_X1 _33266_ (.A(_17101_),
    .B(_16943_),
    .Z(_08320_));
 XOR2_X2 _33267_ (.A(_08241_),
    .B(_06927_),
    .Z(_08321_));
 XNOR2_X1 _33268_ (.A(_07564_),
    .B(_01000_),
    .ZN(_08322_));
 XOR2_X1 _33269_ (.A(_08321_),
    .B(_08322_),
    .Z(_08323_));
 XNOR2_X1 _33270_ (.A(_08323_),
    .B(_07351_),
    .ZN(_08324_));
 MUX2_X1 _33271_ (.A(_08320_),
    .B(_08324_),
    .S(_08300_),
    .Z(_00671_));
 XOR2_X1 _33272_ (.A(_17102_),
    .B(_16944_),
    .Z(_08325_));
 XOR2_X1 _33273_ (.A(_07479_),
    .B(_01001_),
    .Z(_08326_));
 XNOR2_X1 _33274_ (.A(_07109_),
    .B(_08241_),
    .ZN(_08328_));
 XNOR2_X1 _33275_ (.A(_08326_),
    .B(_08328_),
    .ZN(_08329_));
 XNOR2_X1 _33276_ (.A(_07566_),
    .B(_07884_),
    .ZN(_08330_));
 XNOR2_X1 _33277_ (.A(_08329_),
    .B(_08330_),
    .ZN(_08331_));
 MUX2_X1 _33278_ (.A(_08325_),
    .B(_08331_),
    .S(_08300_),
    .Z(_00672_));
 XOR2_X1 _33279_ (.A(_17103_),
    .B(_16945_),
    .Z(_08332_));
 XNOR2_X1 _33280_ (.A(_07702_),
    .B(_01002_),
    .ZN(_08333_));
 XNOR2_X1 _33281_ (.A(_07884_),
    .B(_07628_),
    .ZN(_08334_));
 XNOR2_X1 _33282_ (.A(_08333_),
    .B(_08334_),
    .ZN(_08335_));
 XNOR2_X1 _33283_ (.A(_08335_),
    .B(_08126_),
    .ZN(_08336_));
 MUX2_X1 _33284_ (.A(_08332_),
    .B(_08336_),
    .S(_08300_),
    .Z(_00673_));
 XOR2_X1 _33285_ (.A(_17104_),
    .B(_16947_),
    .Z(_08338_));
 XNOR2_X1 _33286_ (.A(_08296_),
    .B(_15346_),
    .ZN(_08339_));
 XNOR2_X1 _33287_ (.A(_08010_),
    .B(_08339_),
    .ZN(_08340_));
 XOR2_X2 _33288_ (.A(_08125_),
    .B(_07825_),
    .Z(_08341_));
 XNOR2_X1 _33289_ (.A(_08340_),
    .B(_08341_),
    .ZN(_08342_));
 MUX2_X1 _33290_ (.A(_08338_),
    .B(_08342_),
    .S(_08300_),
    .Z(_00674_));
 XOR2_X1 _33291_ (.A(_17105_),
    .B(_16948_),
    .Z(_08343_));
 XNOR2_X1 _33292_ (.A(_08068_),
    .B(_01004_),
    .ZN(_08344_));
 XNOR2_X1 _33293_ (.A(_08185_),
    .B(_08344_),
    .ZN(_08345_));
 XNOR2_X1 _33294_ (.A(_08296_),
    .B(_05983_),
    .ZN(_08347_));
 XNOR2_X1 _33295_ (.A(_08345_),
    .B(_08347_),
    .ZN(_08348_));
 MUX2_X1 _33296_ (.A(_08343_),
    .B(_08348_),
    .S(_08300_),
    .Z(_00675_));
 XOR2_X1 _33297_ (.A(_17106_),
    .B(_16949_),
    .Z(_08349_));
 XOR2_X1 _33298_ (.A(_08309_),
    .B(_01005_),
    .Z(_08350_));
 XNOR2_X1 _33299_ (.A(_05369_),
    .B(_06667_),
    .ZN(_08351_));
 XNOR2_X1 _33300_ (.A(_08351_),
    .B(_08184_),
    .ZN(_08352_));
 XNOR2_X1 _33301_ (.A(_08350_),
    .B(_08352_),
    .ZN(_08353_));
 MUX2_X1 _33302_ (.A(_08349_),
    .B(_08353_),
    .S(_08300_),
    .Z(_00636_));
 XOR2_X1 _33303_ (.A(_17107_),
    .B(_16950_),
    .Z(_08354_));
 XNOR2_X1 _33304_ (.A(_08184_),
    .B(_05734_),
    .ZN(_08356_));
 XNOR2_X1 _33305_ (.A(_06437_),
    .B(_01006_),
    .ZN(_08357_));
 XOR2_X1 _33306_ (.A(_08356_),
    .B(_08357_),
    .Z(_08358_));
 XNOR2_X1 _33307_ (.A(_08315_),
    .B(_08309_),
    .ZN(_08359_));
 XNOR2_X1 _33308_ (.A(_08358_),
    .B(_08359_),
    .ZN(_08360_));
 BUF_X2 _33309_ (.A(_09038_),
    .Z(_08361_));
 MUX2_X1 _33310_ (.A(_08354_),
    .B(_08360_),
    .S(_08361_),
    .Z(_00637_));
 XOR2_X1 _33311_ (.A(_17108_),
    .B(_16951_),
    .Z(_08362_));
 XOR2_X2 _33312_ (.A(_07193_),
    .B(_06927_),
    .Z(_08363_));
 XNOR2_X1 _33313_ (.A(_08363_),
    .B(_06351_),
    .ZN(_08364_));
 XNOR2_X1 _33314_ (.A(_06835_),
    .B(_01007_),
    .ZN(_08366_));
 XNOR2_X1 _33315_ (.A(_08366_),
    .B(_06553_),
    .ZN(_08367_));
 XNOR2_X1 _33316_ (.A(_08364_),
    .B(_08367_),
    .ZN(_08368_));
 MUX2_X1 _33317_ (.A(_08362_),
    .B(_08368_),
    .S(_08361_),
    .Z(_00638_));
 XOR2_X1 _33318_ (.A(_17109_),
    .B(_16952_),
    .Z(_08369_));
 XNOR2_X1 _33319_ (.A(_08184_),
    .B(_06757_),
    .ZN(_08370_));
 XNOR2_X1 _33320_ (.A(_07269_),
    .B(_15912_),
    .ZN(_08371_));
 XNOR2_X1 _33321_ (.A(_08370_),
    .B(_08371_),
    .ZN(_08372_));
 XNOR2_X1 _33322_ (.A(_07109_),
    .B(_07564_),
    .ZN(_08373_));
 XNOR2_X1 _33323_ (.A(_08321_),
    .B(_08373_),
    .ZN(_08374_));
 XNOR2_X1 _33324_ (.A(_08372_),
    .B(_08374_),
    .ZN(_08376_));
 MUX2_X1 _33325_ (.A(_08369_),
    .B(_08376_),
    .S(_08361_),
    .Z(_00639_));
 XOR2_X1 _33326_ (.A(_08184_),
    .B(_07349_),
    .Z(_08377_));
 XNOR2_X1 _33327_ (.A(_08377_),
    .B(_08334_),
    .ZN(_08378_));
 XNOR2_X1 _33328_ (.A(_07478_),
    .B(_01009_),
    .ZN(_08379_));
 XNOR2_X1 _33329_ (.A(_08328_),
    .B(_08379_),
    .ZN(_08380_));
 OR2_X1 _33330_ (.A1(_08378_),
    .A2(_08380_),
    .ZN(_08381_));
 AOI21_X1 _33331_ (.A(_01331_),
    .B1(_08378_),
    .B2(_08380_),
    .ZN(_08382_));
 XNOR2_X1 _33332_ (.A(_17111_),
    .B(_16953_),
    .ZN(_08383_));
 AOI22_X1 _33333_ (.A1(_08381_),
    .A2(_08382_),
    .B1(_01331_),
    .B2(_08383_),
    .ZN(_00640_));
 XOR2_X1 _33334_ (.A(_17112_),
    .B(_16954_),
    .Z(_08385_));
 XNOR2_X1 _33335_ (.A(_08341_),
    .B(_07419_),
    .ZN(_08386_));
 XNOR2_X1 _33336_ (.A(_07628_),
    .B(_01010_),
    .ZN(_08387_));
 XNOR2_X1 _33337_ (.A(_08387_),
    .B(_07756_),
    .ZN(_08388_));
 XNOR2_X1 _33338_ (.A(_08386_),
    .B(_08388_),
    .ZN(_08389_));
 MUX2_X1 _33339_ (.A(_08385_),
    .B(_08389_),
    .S(_08361_),
    .Z(_00641_));
 XOR2_X1 _33340_ (.A(_17113_),
    .B(_16955_),
    .Z(_08390_));
 XNOR2_X1 _33341_ (.A(_07702_),
    .B(_08068_),
    .ZN(_08391_));
 XNOR2_X1 _33342_ (.A(_08391_),
    .B(_08296_),
    .ZN(_08392_));
 XNOR2_X1 _33343_ (.A(_07825_),
    .B(_01011_),
    .ZN(_08393_));
 XOR2_X1 _33344_ (.A(_08393_),
    .B(_07940_),
    .Z(_08395_));
 XNOR2_X1 _33345_ (.A(_08392_),
    .B(_08395_),
    .ZN(_08396_));
 MUX2_X1 _33346_ (.A(_08390_),
    .B(_08396_),
    .S(_08361_),
    .Z(_00642_));
 XOR2_X1 _33347_ (.A(_17114_),
    .B(_16956_),
    .Z(_08397_));
 XNOR2_X1 _33348_ (.A(_08068_),
    .B(_05484_),
    .ZN(_08398_));
 XNOR2_X1 _33349_ (.A(_08398_),
    .B(_08241_),
    .ZN(_08399_));
 XNOR2_X1 _33350_ (.A(_05983_),
    .B(_01012_),
    .ZN(_08400_));
 XNOR2_X1 _33351_ (.A(_08400_),
    .B(_08009_),
    .ZN(_08401_));
 XNOR2_X1 _33352_ (.A(_08399_),
    .B(_08401_),
    .ZN(_08402_));
 MUX2_X1 _33353_ (.A(_08397_),
    .B(_08402_),
    .S(_08361_),
    .Z(_00643_));
 XOR2_X1 _33354_ (.A(_17115_),
    .B(_16958_),
    .Z(_08404_));
 XNOR2_X1 _33355_ (.A(_08185_),
    .B(_05734_),
    .ZN(_08405_));
 XNOR2_X1 _33356_ (.A(_08405_),
    .B(_06233_),
    .ZN(_08406_));
 XNOR2_X1 _33357_ (.A(_08406_),
    .B(_06667_),
    .ZN(_08407_));
 XNOR2_X1 _33358_ (.A(_08407_),
    .B(_01014_),
    .ZN(_08408_));
 MUX2_X1 _33359_ (.A(_08404_),
    .B(_08408_),
    .S(_08361_),
    .Z(_00604_));
 XOR2_X1 _33360_ (.A(_17116_),
    .B(_16959_),
    .Z(_08409_));
 XOR2_X1 _33361_ (.A(_08315_),
    .B(_06351_),
    .Z(_08410_));
 XNOR2_X1 _33362_ (.A(_05485_),
    .B(_08356_),
    .ZN(_08411_));
 XNOR2_X1 _33363_ (.A(_08410_),
    .B(_08411_),
    .ZN(_08412_));
 INV_X1 _33364_ (.A(_01016_),
    .ZN(_08414_));
 XNOR2_X1 _33365_ (.A(_08412_),
    .B(_08414_),
    .ZN(_08415_));
 MUX2_X1 _33366_ (.A(_08409_),
    .B(_08415_),
    .S(_08361_),
    .Z(_00605_));
 XOR2_X1 _33367_ (.A(_17117_),
    .B(_16960_),
    .Z(_08416_));
 XNOR2_X1 _33368_ (.A(_06438_),
    .B(_01018_),
    .ZN(_08417_));
 XNOR2_X1 _33369_ (.A(_08363_),
    .B(_06757_),
    .ZN(_08418_));
 XNOR2_X1 _33370_ (.A(_08417_),
    .B(_08418_),
    .ZN(_08419_));
 MUX2_X1 _33371_ (.A(_08416_),
    .B(_08419_),
    .S(_08361_),
    .Z(_00606_));
 XOR2_X1 _33372_ (.A(_17118_),
    .B(_16961_),
    .Z(_08420_));
 XNOR2_X1 _33373_ (.A(_07349_),
    .B(_01020_),
    .ZN(_08421_));
 XOR2_X1 _33374_ (.A(_07023_),
    .B(_08421_),
    .Z(_08423_));
 XNOR2_X1 _33375_ (.A(_08370_),
    .B(_08373_),
    .ZN(_08424_));
 XNOR2_X1 _33376_ (.A(_08423_),
    .B(_08424_),
    .ZN(_08425_));
 MUX2_X1 _33377_ (.A(_08420_),
    .B(_08425_),
    .S(_08361_),
    .Z(_00607_));
 XOR2_X1 _33378_ (.A(_17119_),
    .B(_16962_),
    .Z(_08426_));
 XOR2_X1 _33379_ (.A(_07419_),
    .B(_01022_),
    .Z(_08427_));
 XOR2_X1 _33380_ (.A(_07481_),
    .B(_08427_),
    .Z(_08428_));
 XNOR2_X1 _33381_ (.A(_08378_),
    .B(_08428_),
    .ZN(_08429_));
 MUX2_X1 _33382_ (.A(_08426_),
    .B(_08429_),
    .S(_09039_),
    .Z(_00608_));
 XOR2_X1 _33383_ (.A(_17120_),
    .B(_16963_),
    .Z(_08430_));
 XNOR2_X1 _33384_ (.A(_07825_),
    .B(_01024_),
    .ZN(_08432_));
 XNOR2_X1 _33385_ (.A(_08432_),
    .B(_07702_),
    .ZN(_08433_));
 XNOR2_X1 _33386_ (.A(_07479_),
    .B(_08125_),
    .ZN(_08434_));
 XNOR2_X1 _33387_ (.A(_08433_),
    .B(_08434_),
    .ZN(_08435_));
 MUX2_X1 _33388_ (.A(_08430_),
    .B(_08435_),
    .S(_09039_),
    .Z(_00609_));
 XOR2_X1 _33389_ (.A(_17122_),
    .B(_16964_),
    .Z(_08436_));
 XNOR2_X1 _33390_ (.A(_08296_),
    .B(_01026_),
    .ZN(_08437_));
 XNOR2_X1 _33391_ (.A(_07757_),
    .B(_08437_),
    .ZN(_08438_));
 XNOR2_X1 _33392_ (.A(_08068_),
    .B(_08009_),
    .ZN(_08439_));
 XNOR2_X1 _33393_ (.A(_08438_),
    .B(_08439_),
    .ZN(_08440_));
 MUX2_X1 _33394_ (.A(_08436_),
    .B(_08440_),
    .S(_09039_),
    .Z(_00610_));
 XOR2_X1 _33395_ (.A(_17123_),
    .B(_16965_),
    .Z(_08442_));
 XOR2_X1 _33396_ (.A(_08184_),
    .B(_01028_),
    .Z(_08443_));
 XNOR2_X1 _33397_ (.A(_08443_),
    .B(_08010_),
    .ZN(_08444_));
 XNOR2_X1 _33398_ (.A(_08307_),
    .B(_05983_),
    .ZN(_08445_));
 XNOR2_X1 _33399_ (.A(_08444_),
    .B(_08445_),
    .ZN(_08446_));
 MUX2_X1 _33400_ (.A(_08442_),
    .B(_08446_),
    .S(_09039_),
    .Z(_00611_));
 AND3_X1 _33401_ (.A1(_05071_),
    .A2(_05072_),
    .A3(_01198_),
    .ZN(_00603_));
 XNOR2_X1 _33402_ (.A(_05369_),
    .B(_01014_),
    .ZN(_00884_));
 XNOR2_X1 _33403_ (.A(_06437_),
    .B(_08414_),
    .ZN(_00885_));
 XNOR2_X1 _33404_ (.A(_06835_),
    .B(_03639_),
    .ZN(_00886_));
 XOR2_X1 _33405_ (.A(_07269_),
    .B(_17118_),
    .Z(_00887_));
 XNOR2_X1 _33406_ (.A(_07478_),
    .B(_17119_),
    .ZN(_00888_));
 XOR2_X1 _33407_ (.A(_07756_),
    .B(_01024_),
    .Z(_00889_));
 XOR2_X1 _33408_ (.A(_07940_),
    .B(_01026_),
    .Z(_00890_));
 XNOR2_X1 _33409_ (.A(_05484_),
    .B(_17123_),
    .ZN(_00891_));
 XOR2_X1 _33410_ (.A(_02050_),
    .B(_01042_),
    .Z(_00980_));
 XNOR2_X1 _33411_ (.A(_03042_),
    .B(_05042_),
    .ZN(_00981_));
 XNOR2_X1 _33412_ (.A(_03446_),
    .B(_17149_),
    .ZN(_00982_));
 XNOR2_X1 _33413_ (.A(_03821_),
    .B(_01662_),
    .ZN(_00983_));
 XNOR2_X1 _33414_ (.A(_04248_),
    .B(_17151_),
    .ZN(_00984_));
 XOR2_X1 _33415_ (.A(_04385_),
    .B(_01044_),
    .Z(_00985_));
 XOR2_X1 _33416_ (.A(_04562_),
    .B(_01048_),
    .Z(_00986_));
 XNOR2_X1 _33417_ (.A(_02139_),
    .B(_17155_),
    .ZN(_00987_));
 XOR2_X1 _33418_ (.A(_11776_),
    .B(_01033_),
    .Z(_00940_));
 XNOR2_X1 _33419_ (.A(_12181_),
    .B(_01793_),
    .ZN(_00941_));
 XNOR2_X1 _33420_ (.A(_12575_),
    .B(_17181_),
    .ZN(_00942_));
 XNOR2_X1 _33421_ (.A(_12952_),
    .B(_17182_),
    .ZN(_00943_));
 XNOR2_X1 _33422_ (.A(_13159_),
    .B(_17183_),
    .ZN(_00944_));
 XOR2_X1 _33423_ (.A(_13463_),
    .B(_01035_),
    .Z(_00945_));
 XNOR2_X1 _33424_ (.A(_13685_),
    .B(_01036_),
    .ZN(_00946_));
 XNOR2_X1 _33425_ (.A(_11877_),
    .B(_17187_),
    .ZN(_00947_));
 XOR2_X1 _33426_ (.A(_08722_),
    .B(_01054_),
    .Z(_00908_));
 XOR2_X1 _33427_ (.A(_09447_),
    .B(_01055_),
    .Z(_00909_));
 XNOR2_X1 _33428_ (.A(_09603_),
    .B(_17085_),
    .ZN(_00910_));
 XNOR2_X1 _33429_ (.A(_09836_),
    .B(_17086_),
    .ZN(_00911_));
 XNOR2_X1 _33430_ (.A(_10181_),
    .B(_17087_),
    .ZN(_00912_));
 XOR2_X1 _33431_ (.A(_10485_),
    .B(_01056_),
    .Z(_00913_));
 XOR2_X1 _33432_ (.A(_10604_),
    .B(_01057_),
    .Z(_00914_));
 XNOR2_X1 _33433_ (.A(_08811_),
    .B(_17091_),
    .ZN(_00915_));
 XNOR2_X1 _33434_ (.A(_05734_),
    .B(_01005_),
    .ZN(_00876_));
 XNOR2_X1 _33435_ (.A(_06351_),
    .B(_15749_),
    .ZN(_00877_));
 XNOR2_X1 _33436_ (.A(_06757_),
    .B(_17108_),
    .ZN(_00878_));
 XNOR2_X1 _33437_ (.A(_07349_),
    .B(_17109_),
    .ZN(_00879_));
 XNOR2_X1 _33438_ (.A(_07419_),
    .B(_17111_),
    .ZN(_00880_));
 XOR2_X1 _33439_ (.A(_07702_),
    .B(_01010_),
    .Z(_00881_));
 XNOR2_X1 _33440_ (.A(_08009_),
    .B(_16111_),
    .ZN(_00882_));
 XNOR2_X1 _33441_ (.A(_08184_),
    .B(_17114_),
    .ZN(_00883_));
 XNOR2_X1 _33442_ (.A(_02617_),
    .B(_01038_),
    .ZN(_00972_));
 XNOR2_X1 _33443_ (.A(_02963_),
    .B(_04984_),
    .ZN(_00973_));
 XNOR2_X1 _33444_ (.A(_03372_),
    .B(_17140_),
    .ZN(_00974_));
 XNOR2_X1 _33445_ (.A(_03902_),
    .B(_01769_),
    .ZN(_00975_));
 XNOR2_X1 _33446_ (.A(_04184_),
    .B(_17143_),
    .ZN(_00976_));
 XNOR2_X1 _33447_ (.A(_04445_),
    .B(_05014_),
    .ZN(_00977_));
 XOR2_X1 _33448_ (.A(_04622_),
    .B(_01041_),
    .Z(_00978_));
 XNOR2_X1 _33449_ (.A(_04859_),
    .B(_17146_),
    .ZN(_00979_));
 XOR2_X1 _33450_ (.A(_11312_),
    .B(_01029_),
    .Z(_00932_));
 XOR2_X1 _33451_ (.A(_12284_),
    .B(_01030_),
    .Z(_00933_));
 XNOR2_X1 _33452_ (.A(_12650_),
    .B(_17172_),
    .ZN(_00934_));
 XNOR2_X1 _33453_ (.A(_12883_),
    .B(_17173_),
    .ZN(_00935_));
 XNOR2_X1 _33454_ (.A(_13216_),
    .B(_17175_),
    .ZN(_00936_));
 XOR2_X1 _33455_ (.A(_13408_),
    .B(_01031_),
    .Z(_00937_));
 XOR2_X1 _33456_ (.A(_13637_),
    .B(_01032_),
    .Z(_00938_));
 XNOR2_X1 _33457_ (.A(_13895_),
    .B(_17178_),
    .ZN(_00939_));
 XOR2_X1 _33458_ (.A(_08502_),
    .B(_01050_),
    .Z(_00900_));
 XOR2_X1 _33459_ (.A(_09372_),
    .B(_01051_),
    .Z(_00901_));
 XNOR2_X1 _33460_ (.A(_09534_),
    .B(_16188_),
    .ZN(_00902_));
 XNOR2_X1 _33461_ (.A(_09914_),
    .B(_17077_),
    .ZN(_00903_));
 XNOR2_X1 _33462_ (.A(_10237_),
    .B(_17079_),
    .ZN(_00904_));
 XOR2_X1 _33463_ (.A(_10431_),
    .B(_01052_),
    .Z(_00905_));
 XOR2_X1 _33464_ (.A(_10651_),
    .B(_01053_),
    .Z(_00906_));
 XNOR2_X1 _33465_ (.A(_10824_),
    .B(_17082_),
    .ZN(_00907_));
 XNOR2_X1 _33466_ (.A(_06233_),
    .B(_17129_),
    .ZN(_00868_));
 XNOR2_X1 _33467_ (.A(_06553_),
    .B(_17130_),
    .ZN(_00869_));
 XNOR2_X1 _33468_ (.A(_06927_),
    .B(_17100_),
    .ZN(_00870_));
 XNOR2_X1 _33469_ (.A(_07109_),
    .B(_17101_),
    .ZN(_00871_));
 XNOR2_X1 _33470_ (.A(_07628_),
    .B(_17102_),
    .ZN(_00872_));
 XOR2_X1 _33471_ (.A(_07825_),
    .B(_17103_),
    .Z(_00873_));
 XOR2_X1 _33472_ (.A(_08068_),
    .B(_17104_),
    .Z(_00874_));
 XNOR2_X1 _33473_ (.A(_08241_),
    .B(_17105_),
    .ZN(_00875_));
 XNOR2_X1 _33474_ (.A(_02385_),
    .B(_17161_),
    .ZN(_00956_));
 XNOR2_X1 _33475_ (.A(_03139_),
    .B(_17162_),
    .ZN(_00957_));
 XNOR2_X1 _33476_ (.A(_03524_),
    .B(_17132_),
    .ZN(_00958_));
 XNOR2_X1 _33477_ (.A(_03745_),
    .B(_17133_),
    .ZN(_00959_));
 XNOR2_X1 _33478_ (.A(_04046_),
    .B(_17134_),
    .ZN(_00960_));
 XNOR2_X1 _33479_ (.A(_04323_),
    .B(_04962_),
    .ZN(_00961_));
 XNOR2_X1 _33480_ (.A(_04689_),
    .B(_17136_),
    .ZN(_00962_));
 XNOR2_X1 _33481_ (.A(_04805_),
    .B(_17137_),
    .ZN(_00963_));
 XNOR2_X1 _33482_ (.A(_11548_),
    .B(_17193_),
    .ZN(_00924_));
 XNOR2_X1 _33483_ (.A(_12385_),
    .B(_17194_),
    .ZN(_00925_));
 XNOR2_X1 _33484_ (.A(_12727_),
    .B(_17164_),
    .ZN(_00926_));
 XNOR2_X1 _33485_ (.A(_13094_),
    .B(_17165_),
    .ZN(_00927_));
 XNOR2_X1 _33486_ (.A(_13346_),
    .B(_01755_),
    .ZN(_00928_));
 XNOR2_X1 _33487_ (.A(_13580_),
    .B(_17167_),
    .ZN(_00929_));
 XNOR2_X1 _33488_ (.A(_13736_),
    .B(_17168_),
    .ZN(_00930_));
 XNOR2_X1 _33489_ (.A(_13842_),
    .B(_17169_),
    .ZN(_00931_));
 XNOR2_X1 _33490_ (.A(_06677_),
    .B(_10932_),
    .ZN(_00892_));
 XNOR2_X1 _33491_ (.A(_09258_),
    .B(_10938_),
    .ZN(_00893_));
 XNOR2_X1 _33492_ (.A(_09685_),
    .B(_17068_),
    .ZN(_00894_));
 XNOR2_X1 _33493_ (.A(_10060_),
    .B(_17069_),
    .ZN(_00895_));
 XNOR2_X1 _33494_ (.A(_10119_),
    .B(_17070_),
    .ZN(_00896_));
 XNOR2_X1 _33495_ (.A(_10371_),
    .B(_17071_),
    .ZN(_00897_));
 XNOR2_X1 _33496_ (.A(_10705_),
    .B(_17072_),
    .ZN(_00898_));
 XNOR2_X1 _33497_ (.A(_10871_),
    .B(_17073_),
    .ZN(_00899_));
 XNOR2_X1 _33498_ (.A(_06667_),
    .B(_17099_),
    .ZN(_00860_));
 XOR2_X1 _33499_ (.A(_07017_),
    .B(_17110_),
    .Z(_00861_));
 XOR2_X1 _33500_ (.A(_07193_),
    .B(_17121_),
    .Z(_00862_));
 XNOR2_X1 _33501_ (.A(_07564_),
    .B(_17124_),
    .ZN(_00863_));
 XNOR2_X1 _33502_ (.A(_07884_),
    .B(_17125_),
    .ZN(_00864_));
 XOR2_X1 _33503_ (.A(_08125_),
    .B(_17126_),
    .Z(_00865_));
 XNOR2_X1 _33504_ (.A(_08296_),
    .B(_17127_),
    .ZN(_00866_));
 XNOR2_X1 _33505_ (.A(_05983_),
    .B(_17128_),
    .ZN(_00867_));
 XNOR2_X1 _33506_ (.A(_03252_),
    .B(_02839_),
    .ZN(_00948_));
 XOR2_X1 _33507_ (.A(_03615_),
    .B(_17142_),
    .Z(_00949_));
 XNOR2_X1 _33508_ (.A(_03982_),
    .B(_03618_),
    .ZN(_00950_));
 XNOR2_X1 _33509_ (.A(_04112_),
    .B(_17156_),
    .ZN(_00951_));
 XNOR2_X1 _33510_ (.A(_04500_),
    .B(_17157_),
    .ZN(_00952_));
 XOR2_X1 _33511_ (.A(_04745_),
    .B(_17158_),
    .Z(_00953_));
 XNOR2_X1 _33512_ (.A(_04924_),
    .B(_17159_),
    .ZN(_00954_));
 XOR2_X1 _33513_ (.A(_02837_),
    .B(_17160_),
    .Z(_00955_));
 XNOR2_X1 _33514_ (.A(_12499_),
    .B(_17163_),
    .ZN(_00916_));
 XNOR2_X1 _33515_ (.A(_12807_),
    .B(_01730_),
    .ZN(_00917_));
 XNOR2_X1 _33516_ (.A(_13017_),
    .B(_01733_),
    .ZN(_00918_));
 XNOR2_X1 _33517_ (.A(_13287_),
    .B(_17188_),
    .ZN(_00919_));
 XNOR2_X1 _33518_ (.A(_13515_),
    .B(_17189_),
    .ZN(_00920_));
 XNOR2_X1 _33519_ (.A(_13791_),
    .B(_01742_),
    .ZN(_00921_));
 XNOR2_X1 _33520_ (.A(_13946_),
    .B(_13793_),
    .ZN(_00922_));
 XNOR2_X1 _33521_ (.A(_12101_),
    .B(_17192_),
    .ZN(_00923_));
 XNOR2_X1 _33522_ (.A(_09147_),
    .B(_04132_),
    .ZN(_00964_));
 XNOR2_X1 _33523_ (.A(_09758_),
    .B(_09041_),
    .ZN(_00965_));
 XNOR2_X1 _33524_ (.A(_09984_),
    .B(_17089_),
    .ZN(_00966_));
 XNOR2_X1 _33525_ (.A(_10307_),
    .B(_17092_),
    .ZN(_00967_));
 XNOR2_X1 _33526_ (.A(_10542_),
    .B(_17093_),
    .ZN(_00968_));
 XNOR2_X1 _33527_ (.A(_10770_),
    .B(_14663_),
    .ZN(_00969_));
 XNOR2_X1 _33528_ (.A(_10924_),
    .B(_17095_),
    .ZN(_00970_));
 XNOR2_X1 _33529_ (.A(_09035_),
    .B(_17096_),
    .ZN(_00971_));
 BUF_X2 _33530_ (.A(net2),
    .Z(_01330_));
 BUF_X1 _33531_ (.A(\u0.r0.rcnt[0] ),
    .Z(_17063_));
 CLKBUF_X1 _33532_ (.A(\u0.r0.rcnt[1] ),
    .Z(_17064_));
 CLKBUF_X1 _33533_ (.A(\u0.r0.rcnt[2] ),
    .Z(_17065_));
 CLKBUF_X1 _33534_ (.A(\u0.r0.rcnt[3] ),
    .Z(_17066_));
 CLKBUF_X1 _33535_ (.A(_01186_),
    .Z(_00587_));
 CLKBUF_X1 _33536_ (.A(_01187_),
    .Z(_00588_));
 CLKBUF_X1 _33537_ (.A(_01188_),
    .Z(_00589_));
 CLKBUF_X1 _33538_ (.A(_01189_),
    .Z(_00590_));
 CLKBUF_X1 _33539_ (.A(_01190_),
    .Z(_00591_));
 CLKBUF_X1 _33540_ (.A(_01191_),
    .Z(_00592_));
 CLKBUF_X1 _33541_ (.A(_01192_),
    .Z(_00593_));
 CLKBUF_X1 _33542_ (.A(_01193_),
    .Z(_00594_));
 CLKBUF_X1 _33543_ (.A(_01194_),
    .Z(_00595_));
 CLKBUF_X1 _33544_ (.A(_01195_),
    .Z(_00596_));
 CLKBUF_X1 _33545_ (.A(_01196_),
    .Z(_00597_));
 CLKBUF_X1 _33546_ (.A(_01197_),
    .Z(_00598_));
 CLKBUF_X2 _33547_ (.A(\sa03[0] ),
    .Z(_16703_));
 CLKBUF_X1 _33548_ (.A(\sa03[1] ),
    .Z(_16704_));
 CLKBUF_X2 _33549_ (.A(\sa03[3] ),
    .Z(_16706_));
 CLKBUF_X2 _33550_ (.A(\sa03[2] ),
    .Z(_16705_));
 CLKBUF_X1 _33551_ (.A(\sa03[5] ),
    .Z(_16708_));
 CLKBUF_X1 _33552_ (.A(\sa03[4] ),
    .Z(_16707_));
 CLKBUF_X1 _33553_ (.A(\sa03[7] ),
    .Z(_16710_));
 CLKBUF_X1 _33554_ (.A(\sa03[6] ),
    .Z(_16709_));
 CLKBUF_X1 _33555_ (.A(\sa10[5] ),
    .Z(_16716_));
 CLKBUF_X1 _33556_ (.A(\sa10[4] ),
    .Z(_16715_));
 CLKBUF_X1 _33557_ (.A(\sa10[7] ),
    .Z(_16718_));
 CLKBUF_X1 _33558_ (.A(\sa10[6] ),
    .Z(_16717_));
 CLKBUF_X2 _33559_ (.A(\sa10[1] ),
    .Z(_16712_));
 BUF_X1 _33560_ (.A(\sa10[0] ),
    .Z(_16711_));
 CLKBUF_X2 _33561_ (.A(\sa10[2] ),
    .Z(_16713_));
 CLKBUF_X2 _33562_ (.A(\sa10[3] ),
    .Z(_16714_));
 CLKBUF_X1 _33563_ (.A(\sa21[5] ),
    .Z(_16756_));
 CLKBUF_X1 _33564_ (.A(\sa21[4] ),
    .Z(_16755_));
 CLKBUF_X1 _33565_ (.A(\sa21[7] ),
    .Z(_16758_));
 BUF_X1 _33566_ (.A(\sa21[6] ),
    .Z(_16757_));
 CLKBUF_X2 _33567_ (.A(\sa21[1] ),
    .Z(_16752_));
 CLKBUF_X2 _33568_ (.A(\sa21[0] ),
    .Z(_16751_));
 BUF_X1 _33569_ (.A(\sa21[2] ),
    .Z(_16753_));
 CLKBUF_X2 _33570_ (.A(\sa21[3] ),
    .Z(_16754_));
 BUF_X2 _33571_ (.A(\sa32[0] ),
    .Z(_16791_));
 CLKBUF_X2 _33572_ (.A(\sa32[1] ),
    .Z(_16792_));
 BUF_X1 _33573_ (.A(\sa32[3] ),
    .Z(_16794_));
 CLKBUF_X2 _33574_ (.A(\sa32[2] ),
    .Z(_16793_));
 CLKBUF_X1 _33575_ (.A(\sa32[5] ),
    .Z(_16796_));
 CLKBUF_X1 _33576_ (.A(\sa32[4] ),
    .Z(_16795_));
 CLKBUF_X1 _33577_ (.A(\sa32[7] ),
    .Z(_16798_));
 CLKBUF_X1 _33578_ (.A(\sa32[6] ),
    .Z(_16797_));
 BUF_X2 _33579_ (.A(\u0.tmp_w[0] ),
    .Z(_17067_));
 CLKBUF_X1 _33580_ (.A(\text_in_r[0] ),
    .Z(_16935_));
 BUF_X1 _33581_ (.A(ld_r),
    .Z(_01331_));
 CLKBUF_X1 _33582_ (.A(_00724_),
    .Z(_00125_));
 BUF_X2 _33583_ (.A(\u0.tmp_w[1] ),
    .Z(_17078_));
 CLKBUF_X1 _33584_ (.A(\text_in_r[1] ),
    .Z(_16974_));
 CLKBUF_X1 _33585_ (.A(_00725_),
    .Z(_00126_));
 BUF_X2 _33586_ (.A(\u0.tmp_w[2] ),
    .Z(_17089_));
 CLKBUF_X1 _33587_ (.A(\text_in_r[2] ),
    .Z(_16985_));
 CLKBUF_X1 _33588_ (.A(_00726_),
    .Z(_00127_));
 BUF_X2 _33589_ (.A(\u0.tmp_w[3] ),
    .Z(_17092_));
 CLKBUF_X1 _33590_ (.A(\text_in_r[3] ),
    .Z(_16996_));
 CLKBUF_X1 _33591_ (.A(_00727_),
    .Z(_00128_));
 BUF_X2 _33592_ (.A(\u0.tmp_w[4] ),
    .Z(_17093_));
 CLKBUF_X1 _33593_ (.A(\text_in_r[4] ),
    .Z(_17007_));
 CLKBUF_X1 _33594_ (.A(_00728_),
    .Z(_00129_));
 CLKBUF_X2 _33595_ (.A(\u0.tmp_w[5] ),
    .Z(_17094_));
 CLKBUF_X1 _33596_ (.A(\text_in_r[5] ),
    .Z(_17018_));
 CLKBUF_X1 _33597_ (.A(_00729_),
    .Z(_00130_));
 CLKBUF_X2 _33598_ (.A(\u0.tmp_w[6] ),
    .Z(_17095_));
 CLKBUF_X1 _33599_ (.A(\text_in_r[6] ),
    .Z(_17029_));
 CLKBUF_X1 _33600_ (.A(_00730_),
    .Z(_00131_));
 CLKBUF_X2 _33601_ (.A(\u0.tmp_w[7] ),
    .Z(_17096_));
 CLKBUF_X1 _33602_ (.A(\text_in_r[7] ),
    .Z(_17040_));
 CLKBUF_X1 _33603_ (.A(_00731_),
    .Z(_00132_));
 CLKBUF_X1 _33604_ (.A(_00450_),
    .Z(_01049_));
 CLKBUF_X1 _33605_ (.A(\text_in_r[8] ),
    .Z(_17051_));
 CLKBUF_X1 _33606_ (.A(\u0.tmp_w[8] ),
    .Z(_17097_));
 CLKBUF_X1 _33607_ (.A(_00692_),
    .Z(_00093_));
 CLKBUF_X2 _33608_ (.A(\u0.tmp_w[9] ),
    .Z(_17098_));
 CLKBUF_X1 _33609_ (.A(\text_in_r[9] ),
    .Z(_17062_));
 CLKBUF_X1 _33610_ (.A(_00693_),
    .Z(_00094_));
 BUF_X2 _33611_ (.A(\u0.tmp_w[10] ),
    .Z(_17068_));
 CLKBUF_X1 _33612_ (.A(\text_in_r[10] ),
    .Z(_16946_));
 CLKBUF_X1 _33613_ (.A(_00694_),
    .Z(_00095_));
 BUF_X2 _33614_ (.A(\u0.tmp_w[11] ),
    .Z(_17069_));
 CLKBUF_X1 _33615_ (.A(\text_in_r[11] ),
    .Z(_16957_));
 CLKBUF_X1 _33616_ (.A(_00695_),
    .Z(_00096_));
 CLKBUF_X2 _33617_ (.A(\u0.tmp_w[12] ),
    .Z(_17070_));
 CLKBUF_X1 _33618_ (.A(\text_in_r[12] ),
    .Z(_16966_));
 CLKBUF_X1 _33619_ (.A(_00696_),
    .Z(_00097_));
 BUF_X2 _33620_ (.A(\u0.tmp_w[13] ),
    .Z(_17071_));
 CLKBUF_X1 _33621_ (.A(\text_in_r[13] ),
    .Z(_16967_));
 CLKBUF_X1 _33622_ (.A(_00697_),
    .Z(_00098_));
 CLKBUF_X2 _33623_ (.A(\u0.tmp_w[14] ),
    .Z(_17072_));
 CLKBUF_X1 _33624_ (.A(\text_in_r[14] ),
    .Z(_16968_));
 CLKBUF_X1 _33625_ (.A(_00698_),
    .Z(_00099_));
 CLKBUF_X2 _33626_ (.A(\u0.tmp_w[15] ),
    .Z(_17073_));
 CLKBUF_X1 _33627_ (.A(\text_in_r[15] ),
    .Z(_16969_));
 CLKBUF_X1 _33628_ (.A(_00699_),
    .Z(_00100_));
 CLKBUF_X1 _33629_ (.A(_00451_),
    .Z(_01050_));
 CLKBUF_X1 _33630_ (.A(\text_in_r[16] ),
    .Z(_16970_));
 CLKBUF_X2 _33631_ (.A(\u0.tmp_w[16] ),
    .Z(_17074_));
 CLKBUF_X1 _33632_ (.A(_00660_),
    .Z(_00061_));
 CLKBUF_X1 _33633_ (.A(_00452_),
    .Z(_01051_));
 CLKBUF_X1 _33634_ (.A(\text_in_r[17] ),
    .Z(_16971_));
 BUF_X2 _33635_ (.A(\u0.tmp_w[17] ),
    .Z(_17075_));
 CLKBUF_X1 _33636_ (.A(_00661_),
    .Z(_00062_));
 BUF_X2 _33637_ (.A(\u0.tmp_w[18] ),
    .Z(_17076_));
 CLKBUF_X1 _33638_ (.A(\text_in_r[18] ),
    .Z(_16972_));
 CLKBUF_X1 _33639_ (.A(_00662_),
    .Z(_00063_));
 BUF_X2 _33640_ (.A(\u0.tmp_w[19] ),
    .Z(_17077_));
 CLKBUF_X1 _33641_ (.A(\text_in_r[19] ),
    .Z(_16973_));
 CLKBUF_X1 _33642_ (.A(_00663_),
    .Z(_00064_));
 CLKBUF_X2 _33643_ (.A(\u0.tmp_w[20] ),
    .Z(_17079_));
 CLKBUF_X1 _33644_ (.A(\text_in_r[20] ),
    .Z(_16975_));
 CLKBUF_X1 _33645_ (.A(_00664_),
    .Z(_00065_));
 CLKBUF_X1 _33646_ (.A(_00453_),
    .Z(_01052_));
 CLKBUF_X1 _33647_ (.A(\text_in_r[21] ),
    .Z(_16976_));
 BUF_X1 _33648_ (.A(\u0.tmp_w[21] ),
    .Z(_17080_));
 CLKBUF_X1 _33649_ (.A(_00665_),
    .Z(_00066_));
 CLKBUF_X1 _33650_ (.A(_00454_),
    .Z(_01053_));
 CLKBUF_X1 _33651_ (.A(\text_in_r[22] ),
    .Z(_16977_));
 BUF_X1 _33652_ (.A(\u0.tmp_w[22] ),
    .Z(_17081_));
 CLKBUF_X1 _33653_ (.A(_00666_),
    .Z(_00067_));
 BUF_X2 _33654_ (.A(\u0.tmp_w[23] ),
    .Z(_17082_));
 CLKBUF_X1 _33655_ (.A(\text_in_r[23] ),
    .Z(_16978_));
 CLKBUF_X1 _33656_ (.A(_00667_),
    .Z(_00068_));
 CLKBUF_X1 _33657_ (.A(_00455_),
    .Z(_01054_));
 CLKBUF_X1 _33658_ (.A(\text_in_r[24] ),
    .Z(_16979_));
 CLKBUF_X2 _33659_ (.A(\u0.tmp_w[24] ),
    .Z(_17083_));
 CLKBUF_X1 _33660_ (.A(_00628_),
    .Z(_00029_));
 CLKBUF_X1 _33661_ (.A(_00456_),
    .Z(_01055_));
 CLKBUF_X1 _33662_ (.A(\text_in_r[25] ),
    .Z(_16980_));
 BUF_X1 _33663_ (.A(\u0.tmp_w[25] ),
    .Z(_17084_));
 CLKBUF_X1 _33664_ (.A(_00629_),
    .Z(_00030_));
 BUF_X2 _33665_ (.A(\u0.tmp_w[26] ),
    .Z(_17085_));
 CLKBUF_X1 _33666_ (.A(\text_in_r[26] ),
    .Z(_16981_));
 CLKBUF_X1 _33667_ (.A(_00630_),
    .Z(_00031_));
 BUF_X2 _33668_ (.A(\u0.tmp_w[27] ),
    .Z(_17086_));
 CLKBUF_X1 _33669_ (.A(\text_in_r[27] ),
    .Z(_16982_));
 CLKBUF_X1 _33670_ (.A(_00631_),
    .Z(_00032_));
 BUF_X2 _33671_ (.A(\u0.tmp_w[28] ),
    .Z(_17087_));
 CLKBUF_X1 _33672_ (.A(\text_in_r[28] ),
    .Z(_16983_));
 CLKBUF_X1 _33673_ (.A(_00632_),
    .Z(_00033_));
 CLKBUF_X1 _33674_ (.A(_00457_),
    .Z(_01056_));
 CLKBUF_X1 _33675_ (.A(\text_in_r[29] ),
    .Z(_16984_));
 BUF_X1 _33676_ (.A(\u0.tmp_w[29] ),
    .Z(_17088_));
 CLKBUF_X1 _33677_ (.A(_00633_),
    .Z(_00034_));
 CLKBUF_X1 _33678_ (.A(_00458_),
    .Z(_01057_));
 CLKBUF_X1 _33679_ (.A(\text_in_r[30] ),
    .Z(_16986_));
 CLKBUF_X2 _33680_ (.A(\u0.tmp_w[30] ),
    .Z(_17090_));
 CLKBUF_X1 _33681_ (.A(_00634_),
    .Z(_00035_));
 BUF_X2 _33682_ (.A(\u0.tmp_w[31] ),
    .Z(_17091_));
 CLKBUF_X1 _33683_ (.A(\text_in_r[31] ),
    .Z(_16987_));
 CLKBUF_X1 _33684_ (.A(_00635_),
    .Z(_00036_));
 CLKBUF_X2 _33685_ (.A(\sa02[0] ),
    .Z(_16695_));
 BUF_X2 _33686_ (.A(\sa02[1] ),
    .Z(_16696_));
 BUF_X2 _33687_ (.A(\sa02[3] ),
    .Z(_16698_));
 CLKBUF_X2 _33688_ (.A(\sa02[2] ),
    .Z(_16697_));
 CLKBUF_X1 _33689_ (.A(\sa02[5] ),
    .Z(_16700_));
 CLKBUF_X1 _33690_ (.A(\sa02[4] ),
    .Z(_16699_));
 CLKBUF_X1 _33691_ (.A(\sa02[7] ),
    .Z(_16702_));
 CLKBUF_X1 _33692_ (.A(\sa02[6] ),
    .Z(_16701_));
 CLKBUF_X1 _33693_ (.A(\sa13[5] ),
    .Z(_16740_));
 CLKBUF_X1 _33694_ (.A(\sa13[4] ),
    .Z(_16739_));
 CLKBUF_X1 _33695_ (.A(\sa13[7] ),
    .Z(_16742_));
 CLKBUF_X1 _33696_ (.A(\sa13[6] ),
    .Z(_16741_));
 CLKBUF_X2 _33697_ (.A(\sa13[1] ),
    .Z(_16736_));
 CLKBUF_X2 _33698_ (.A(\sa13[0] ),
    .Z(_16735_));
 CLKBUF_X2 _33699_ (.A(\sa13[2] ),
    .Z(_16737_));
 CLKBUF_X2 _33700_ (.A(\sa13[3] ),
    .Z(_16738_));
 CLKBUF_X1 _33701_ (.A(\sa20[5] ),
    .Z(_16748_));
 CLKBUF_X1 _33702_ (.A(\sa20[4] ),
    .Z(_16747_));
 BUF_X1 _33703_ (.A(\sa20[7] ),
    .Z(_16750_));
 CLKBUF_X1 _33704_ (.A(\sa20[6] ),
    .Z(_16749_));
 CLKBUF_X2 _33705_ (.A(\sa20[1] ),
    .Z(_16744_));
 CLKBUF_X2 _33706_ (.A(\sa20[0] ),
    .Z(_16743_));
 CLKBUF_X2 _33707_ (.A(\sa20[2] ),
    .Z(_16745_));
 CLKBUF_X2 _33708_ (.A(\sa20[3] ),
    .Z(_16746_));
 CLKBUF_X1 _33709_ (.A(\sa31[0] ),
    .Z(_16783_));
 CLKBUF_X2 _33710_ (.A(\sa31[1] ),
    .Z(_16784_));
 CLKBUF_X2 _33711_ (.A(\sa31[3] ),
    .Z(_16786_));
 CLKBUF_X2 _33712_ (.A(\sa31[2] ),
    .Z(_16785_));
 CLKBUF_X1 _33713_ (.A(\sa31[5] ),
    .Z(_16788_));
 CLKBUF_X1 _33714_ (.A(\sa31[4] ),
    .Z(_16787_));
 BUF_X1 _33715_ (.A(\sa31[7] ),
    .Z(_16790_));
 CLKBUF_X1 _33716_ (.A(\sa31[6] ),
    .Z(_16789_));
 CLKBUF_X2 _33717_ (.A(\u0.w[2][0] ),
    .Z(_17163_));
 CLKBUF_X1 _33718_ (.A(\text_in_r[32] ),
    .Z(_16988_));
 CLKBUF_X1 _33719_ (.A(_00716_),
    .Z(_00117_));
 BUF_X1 _33720_ (.A(\u0.w[2][1] ),
    .Z(_17174_));
 CLKBUF_X1 _33721_ (.A(\text_in_r[33] ),
    .Z(_16989_));
 CLKBUF_X1 _33722_ (.A(_00717_),
    .Z(_00118_));
 BUF_X1 _33723_ (.A(\u0.w[2][2] ),
    .Z(_17185_));
 CLKBUF_X1 _33724_ (.A(\text_in_r[34] ),
    .Z(_16990_));
 CLKBUF_X1 _33725_ (.A(_00718_),
    .Z(_00119_));
 CLKBUF_X2 _33726_ (.A(\u0.w[2][3] ),
    .Z(_17188_));
 CLKBUF_X1 _33727_ (.A(\text_in_r[35] ),
    .Z(_16991_));
 CLKBUF_X1 _33728_ (.A(_00719_),
    .Z(_00120_));
 CLKBUF_X2 _33729_ (.A(\u0.w[2][4] ),
    .Z(_17189_));
 CLKBUF_X1 _33730_ (.A(\text_in_r[36] ),
    .Z(_16992_));
 CLKBUF_X1 _33731_ (.A(_00720_),
    .Z(_00121_));
 BUF_X1 _33732_ (.A(\u0.w[2][5] ),
    .Z(_17190_));
 CLKBUF_X1 _33733_ (.A(\text_in_r[37] ),
    .Z(_16993_));
 CLKBUF_X1 _33734_ (.A(_00721_),
    .Z(_00122_));
 BUF_X1 _33735_ (.A(\u0.w[2][6] ),
    .Z(_17191_));
 CLKBUF_X1 _33736_ (.A(\text_in_r[38] ),
    .Z(_16994_));
 CLKBUF_X1 _33737_ (.A(_00722_),
    .Z(_00123_));
 CLKBUF_X2 _33738_ (.A(\u0.w[2][7] ),
    .Z(_17192_));
 CLKBUF_X1 _33739_ (.A(\text_in_r[39] ),
    .Z(_16995_));
 CLKBUF_X1 _33740_ (.A(_00723_),
    .Z(_00124_));
 CLKBUF_X1 _33741_ (.A(_00389_),
    .Z(_00988_));
 CLKBUF_X1 _33742_ (.A(net34),
    .Z(_01325_));
 CLKBUF_X1 _33743_ (.A(_01058_),
    .Z(_00459_));
 CLKBUF_X1 _33744_ (.A(_00390_),
    .Z(_00989_));
 CLKBUF_X1 _33745_ (.A(net33),
    .Z(_01326_));
 CLKBUF_X1 _33746_ (.A(_01069_),
    .Z(_00470_));
 CLKBUF_X1 _33747_ (.A(_00391_),
    .Z(_00990_));
 BUF_X1 _33748_ (.A(\u0.w[2][8] ),
    .Z(_17193_));
 CLKBUF_X1 _33749_ (.A(\text_in_r[40] ),
    .Z(_16997_));
 CLKBUF_X1 _33750_ (.A(_00684_),
    .Z(_00085_));
 CLKBUF_X1 _33751_ (.A(_00392_),
    .Z(_00991_));
 CLKBUF_X1 _33752_ (.A(net32),
    .Z(_01327_));
 CLKBUF_X1 _33753_ (.A(_01080_),
    .Z(_00481_));
 CLKBUF_X1 _33754_ (.A(_00393_),
    .Z(_00992_));
 CLKBUF_X1 _33755_ (.A(net31),
    .Z(_01328_));
 CLKBUF_X1 _33756_ (.A(_01083_),
    .Z(_00484_));
 CLKBUF_X1 _33757_ (.A(_00394_),
    .Z(_00993_));
 CLKBUF_X1 _33758_ (.A(net30),
    .Z(_01203_));
 CLKBUF_X1 _33759_ (.A(_01084_),
    .Z(_00485_));
 CLKBUF_X1 _33760_ (.A(_00395_),
    .Z(_00994_));
 CLKBUF_X1 _33761_ (.A(net29),
    .Z(_01204_));
 CLKBUF_X1 _33762_ (.A(_01085_),
    .Z(_00486_));
 CLKBUF_X1 _33763_ (.A(_00396_),
    .Z(_00995_));
 CLKBUF_X1 _33764_ (.A(net28),
    .Z(_01205_));
 CLKBUF_X1 _33765_ (.A(_01086_),
    .Z(_00487_));
 CLKBUF_X1 _33766_ (.A(_00397_),
    .Z(_00996_));
 CLKBUF_X1 _33767_ (.A(net27),
    .Z(_01206_));
 CLKBUF_X1 _33768_ (.A(_01087_),
    .Z(_00488_));
 CLKBUF_X1 _33769_ (.A(_00398_),
    .Z(_00997_));
 CLKBUF_X1 _33770_ (.A(net26),
    .Z(_01207_));
 CLKBUF_X1 _33771_ (.A(_01088_),
    .Z(_00489_));
 CLKBUF_X1 _33772_ (.A(_00399_),
    .Z(_00998_));
 CLKBUF_X1 _33773_ (.A(net25),
    .Z(_01208_));
 CLKBUF_X1 _33774_ (.A(_01089_),
    .Z(_00490_));
 CLKBUF_X1 _33775_ (.A(_00400_),
    .Z(_00999_));
 CLKBUF_X1 _33776_ (.A(net24),
    .Z(_01209_));
 CLKBUF_X1 _33777_ (.A(_01059_),
    .Z(_00460_));
 CLKBUF_X1 _33778_ (.A(_00401_),
    .Z(_01000_));
 CLKBUF_X1 _33779_ (.A(net23),
    .Z(_01210_));
 CLKBUF_X1 _33780_ (.A(_01060_),
    .Z(_00461_));
 BUF_X1 _33781_ (.A(\u0.w[2][9] ),
    .Z(_17194_));
 CLKBUF_X1 _33782_ (.A(\text_in_r[41] ),
    .Z(_16998_));
 CLKBUF_X1 _33783_ (.A(_00685_),
    .Z(_00086_));
 CLKBUF_X1 _33784_ (.A(_00402_),
    .Z(_01001_));
 CLKBUF_X1 _33785_ (.A(net22),
    .Z(_01211_));
 CLKBUF_X1 _33786_ (.A(_01061_),
    .Z(_00462_));
 CLKBUF_X1 _33787_ (.A(_00403_),
    .Z(_01002_));
 CLKBUF_X1 _33788_ (.A(net21),
    .Z(_01212_));
 CLKBUF_X1 _33789_ (.A(_01062_),
    .Z(_00463_));
 CLKBUF_X1 _33790_ (.A(_00404_),
    .Z(_01003_));
 CLKBUF_X1 _33791_ (.A(net20),
    .Z(_01214_));
 CLKBUF_X1 _33792_ (.A(_01063_),
    .Z(_00464_));
 CLKBUF_X1 _33793_ (.A(_00405_),
    .Z(_01004_));
 CLKBUF_X1 _33794_ (.A(net19),
    .Z(_01215_));
 CLKBUF_X1 _33795_ (.A(_01064_),
    .Z(_00465_));
 CLKBUF_X1 _33796_ (.A(_00406_),
    .Z(_01005_));
 CLKBUF_X1 _33797_ (.A(net18),
    .Z(_01216_));
 CLKBUF_X1 _33798_ (.A(_01065_),
    .Z(_00466_));
 CLKBUF_X1 _33799_ (.A(_00407_),
    .Z(_01006_));
 CLKBUF_X1 _33800_ (.A(net17),
    .Z(_01217_));
 CLKBUF_X1 _33801_ (.A(_01066_),
    .Z(_00467_));
 CLKBUF_X1 _33802_ (.A(_00408_),
    .Z(_01007_));
 CLKBUF_X1 _33803_ (.A(net16),
    .Z(_01218_));
 CLKBUF_X1 _33804_ (.A(_01067_),
    .Z(_00468_));
 CLKBUF_X1 _33805_ (.A(_00409_),
    .Z(_01008_));
 CLKBUF_X1 _33806_ (.A(net15),
    .Z(_01219_));
 CLKBUF_X1 _33807_ (.A(_01068_),
    .Z(_00469_));
 CLKBUF_X1 _33808_ (.A(_00410_),
    .Z(_01009_));
 CLKBUF_X1 _33809_ (.A(net14),
    .Z(_01220_));
 CLKBUF_X1 _33810_ (.A(_01070_),
    .Z(_00471_));
 CLKBUF_X1 _33811_ (.A(_00411_),
    .Z(_01010_));
 CLKBUF_X1 _33812_ (.A(net13),
    .Z(_01221_));
 CLKBUF_X1 _33813_ (.A(_01071_),
    .Z(_00472_));
 CLKBUF_X2 _33814_ (.A(\u0.w[2][10] ),
    .Z(_17164_));
 CLKBUF_X1 _33815_ (.A(\text_in_r[42] ),
    .Z(_16999_));
 CLKBUF_X1 _33816_ (.A(_00686_),
    .Z(_00087_));
 CLKBUF_X1 _33817_ (.A(_00412_),
    .Z(_01011_));
 CLKBUF_X1 _33818_ (.A(net12),
    .Z(_01222_));
 CLKBUF_X1 _33819_ (.A(_01072_),
    .Z(_00473_));
 CLKBUF_X1 _33820_ (.A(_00413_),
    .Z(_01012_));
 CLKBUF_X1 _33821_ (.A(net11),
    .Z(_01223_));
 CLKBUF_X1 _33822_ (.A(_01073_),
    .Z(_00474_));
 CLKBUF_X1 _33823_ (.A(_00415_),
    .Z(_01014_));
 CLKBUF_X1 _33824_ (.A(_00414_),
    .Z(_01013_));
 CLKBUF_X1 _33825_ (.A(net10),
    .Z(_01225_));
 CLKBUF_X1 _33826_ (.A(_01074_),
    .Z(_00475_));
 CLKBUF_X1 _33827_ (.A(_00417_),
    .Z(_01016_));
 CLKBUF_X1 _33828_ (.A(_00416_),
    .Z(_01015_));
 CLKBUF_X1 _33829_ (.A(net9),
    .Z(_01226_));
 CLKBUF_X1 _33830_ (.A(_01075_),
    .Z(_00476_));
 CLKBUF_X1 _33831_ (.A(_00419_),
    .Z(_01018_));
 CLKBUF_X1 _33832_ (.A(_00418_),
    .Z(_01017_));
 CLKBUF_X1 _33833_ (.A(net8),
    .Z(_01227_));
 CLKBUF_X1 _33834_ (.A(_01076_),
    .Z(_00477_));
 CLKBUF_X1 _33835_ (.A(_00421_),
    .Z(_01020_));
 CLKBUF_X1 _33836_ (.A(_00420_),
    .Z(_01019_));
 CLKBUF_X1 _33837_ (.A(net7),
    .Z(_01228_));
 CLKBUF_X1 _33838_ (.A(_01077_),
    .Z(_00478_));
 CLKBUF_X1 _33839_ (.A(_00423_),
    .Z(_01022_));
 CLKBUF_X1 _33840_ (.A(_00422_),
    .Z(_01021_));
 CLKBUF_X1 _33841_ (.A(net6),
    .Z(_01229_));
 CLKBUF_X1 _33842_ (.A(_01078_),
    .Z(_00479_));
 CLKBUF_X1 _33843_ (.A(_00425_),
    .Z(_01024_));
 CLKBUF_X1 _33844_ (.A(_00424_),
    .Z(_01023_));
 CLKBUF_X1 _33845_ (.A(net5),
    .Z(_01230_));
 CLKBUF_X1 _33846_ (.A(_01079_),
    .Z(_00480_));
 CLKBUF_X1 _33847_ (.A(_00427_),
    .Z(_01026_));
 CLKBUF_X1 _33848_ (.A(_00426_),
    .Z(_01025_));
 CLKBUF_X1 _33849_ (.A(net4),
    .Z(_01231_));
 CLKBUF_X1 _33850_ (.A(_01081_),
    .Z(_00482_));
 CLKBUF_X1 _33851_ (.A(_00429_),
    .Z(_01028_));
 CLKBUF_X1 _33852_ (.A(_00428_),
    .Z(_01027_));
 CLKBUF_X1 _33853_ (.A(net3),
    .Z(_01232_));
 CLKBUF_X1 _33854_ (.A(_01082_),
    .Z(_00483_));
 CLKBUF_X2 _33855_ (.A(\u0.w[2][11] ),
    .Z(_17165_));
 CLKBUF_X1 _33856_ (.A(\text_in_r[43] ),
    .Z(_17000_));
 CLKBUF_X1 _33857_ (.A(_00687_),
    .Z(_00088_));
 BUF_X1 _33858_ (.A(\u0.w[2][12] ),
    .Z(_17166_));
 CLKBUF_X1 _33859_ (.A(\text_in_r[44] ),
    .Z(_17001_));
 CLKBUF_X1 _33860_ (.A(_00688_),
    .Z(_00089_));
 CLKBUF_X2 _33861_ (.A(\u0.w[2][13] ),
    .Z(_17167_));
 CLKBUF_X1 _33862_ (.A(\text_in_r[45] ),
    .Z(_17002_));
 CLKBUF_X1 _33863_ (.A(_00689_),
    .Z(_00090_));
 CLKBUF_X2 _33864_ (.A(\u0.w[2][14] ),
    .Z(_17168_));
 CLKBUF_X1 _33865_ (.A(\text_in_r[46] ),
    .Z(_17003_));
 CLKBUF_X1 _33866_ (.A(_00690_),
    .Z(_00091_));
 CLKBUF_X2 _33867_ (.A(\u0.w[2][15] ),
    .Z(_17169_));
 CLKBUF_X1 _33868_ (.A(\text_in_r[47] ),
    .Z(_17004_));
 CLKBUF_X1 _33869_ (.A(_00691_),
    .Z(_00092_));
 BUF_X1 _33870_ (.A(\u0.w[1][0] ),
    .Z(_17131_));
 BUF_X1 _33871_ (.A(\u0.w[0][0] ),
    .Z(_17099_));
 CLKBUF_X1 _33872_ (.A(net66),
    .Z(_01290_));
 CLKBUF_X1 _33873_ (.A(_01090_),
    .Z(_00491_));
 BUF_X1 _33874_ (.A(\u0.w[1][1] ),
    .Z(_17142_));
 CLKBUF_X1 _33875_ (.A(\u0.w[0][1] ),
    .Z(_17110_));
 CLKBUF_X1 _33876_ (.A(net65),
    .Z(_01291_));
 CLKBUF_X1 _33877_ (.A(_01101_),
    .Z(_00502_));
 BUF_X1 _33878_ (.A(\u0.w[1][2] ),
    .Z(_17153_));
 BUF_X1 _33879_ (.A(\u0.w[0][2] ),
    .Z(_17121_));
 CLKBUF_X1 _33880_ (.A(net64),
    .Z(_01292_));
 CLKBUF_X1 _33881_ (.A(_01112_),
    .Z(_00513_));
 CLKBUF_X2 _33882_ (.A(\u0.w[1][3] ),
    .Z(_17156_));
 BUF_X1 _33883_ (.A(\u0.w[0][3] ),
    .Z(_17124_));
 CLKBUF_X1 _33884_ (.A(net63),
    .Z(_01293_));
 CLKBUF_X1 _33885_ (.A(_01115_),
    .Z(_00516_));
 CLKBUF_X2 _33886_ (.A(\u0.w[1][4] ),
    .Z(_17157_));
 BUF_X1 _33887_ (.A(\u0.w[0][4] ),
    .Z(_17125_));
 CLKBUF_X1 _33888_ (.A(net62),
    .Z(_01294_));
 CLKBUF_X1 _33889_ (.A(_01116_),
    .Z(_00517_));
 CLKBUF_X2 _33890_ (.A(\u0.w[1][5] ),
    .Z(_17158_));
 BUF_X1 _33891_ (.A(\u0.w[0][5] ),
    .Z(_17126_));
 CLKBUF_X1 _33892_ (.A(net61),
    .Z(_01295_));
 CLKBUF_X1 _33893_ (.A(_01117_),
    .Z(_00518_));
 CLKBUF_X2 _33894_ (.A(\u0.w[1][6] ),
    .Z(_17159_));
 BUF_X1 _33895_ (.A(\u0.w[0][6] ),
    .Z(_17127_));
 CLKBUF_X1 _33896_ (.A(net60),
    .Z(_01297_));
 CLKBUF_X1 _33897_ (.A(_01118_),
    .Z(_00519_));
 CLKBUF_X2 _33898_ (.A(\u0.w[1][7] ),
    .Z(_17160_));
 BUF_X1 _33899_ (.A(\u0.w[0][7] ),
    .Z(_17128_));
 CLKBUF_X1 _33900_ (.A(net59),
    .Z(_01298_));
 CLKBUF_X1 _33901_ (.A(_01119_),
    .Z(_00520_));
 BUF_X1 _33902_ (.A(\u0.w[1][8] ),
    .Z(_17161_));
 BUF_X1 _33903_ (.A(\u0.w[0][8] ),
    .Z(_17129_));
 CLKBUF_X1 _33904_ (.A(net58),
    .Z(_01299_));
 CLKBUF_X1 _33905_ (.A(_01120_),
    .Z(_00521_));
 BUF_X1 _33906_ (.A(\u0.w[1][9] ),
    .Z(_17162_));
 CLKBUF_X1 _33907_ (.A(\u0.w[0][9] ),
    .Z(_17130_));
 CLKBUF_X1 _33908_ (.A(net57),
    .Z(_01300_));
 CLKBUF_X1 _33909_ (.A(_01121_),
    .Z(_00522_));
 CLKBUF_X2 _33910_ (.A(\u0.w[1][10] ),
    .Z(_17132_));
 BUF_X1 _33911_ (.A(\u0.w[0][10] ),
    .Z(_17100_));
 CLKBUF_X1 _33912_ (.A(net56),
    .Z(_01301_));
 CLKBUF_X1 _33913_ (.A(_01091_),
    .Z(_00492_));
 CLKBUF_X2 _33914_ (.A(\u0.w[1][11] ),
    .Z(_17133_));
 BUF_X1 _33915_ (.A(\u0.w[0][11] ),
    .Z(_17101_));
 CLKBUF_X1 _33916_ (.A(net55),
    .Z(_01302_));
 CLKBUF_X1 _33917_ (.A(_01092_),
    .Z(_00493_));
 CLKBUF_X2 _33918_ (.A(\u0.w[1][12] ),
    .Z(_17134_));
 BUF_X1 _33919_ (.A(\u0.w[0][12] ),
    .Z(_17102_));
 CLKBUF_X1 _33920_ (.A(net54),
    .Z(_01303_));
 CLKBUF_X1 _33921_ (.A(_01093_),
    .Z(_00494_));
 BUF_X1 _33922_ (.A(\u0.w[1][13] ),
    .Z(_17135_));
 BUF_X1 _33923_ (.A(\u0.w[0][13] ),
    .Z(_17103_));
 CLKBUF_X1 _33924_ (.A(net53),
    .Z(_01304_));
 CLKBUF_X1 _33925_ (.A(_01094_),
    .Z(_00495_));
 CLKBUF_X2 _33926_ (.A(\u0.w[1][14] ),
    .Z(_17136_));
 BUF_X1 _33927_ (.A(\u0.w[0][14] ),
    .Z(_17104_));
 CLKBUF_X1 _33928_ (.A(net52),
    .Z(_01305_));
 CLKBUF_X1 _33929_ (.A(_01095_),
    .Z(_00496_));
 CLKBUF_X2 _33930_ (.A(\u0.w[1][15] ),
    .Z(_17137_));
 BUF_X1 _33931_ (.A(\u0.w[0][15] ),
    .Z(_17105_));
 CLKBUF_X1 _33932_ (.A(net51),
    .Z(_01306_));
 CLKBUF_X1 _33933_ (.A(_01096_),
    .Z(_00497_));
 BUF_X1 _33934_ (.A(\u0.w[1][16] ),
    .Z(_17138_));
 BUF_X1 _33935_ (.A(\u0.w[0][16] ),
    .Z(_17106_));
 CLKBUF_X1 _33936_ (.A(net50),
    .Z(_01308_));
 CLKBUF_X1 _33937_ (.A(_01097_),
    .Z(_00498_));
 CLKBUF_X1 _33938_ (.A(\u0.w[1][17] ),
    .Z(_17139_));
 CLKBUF_X1 _33939_ (.A(\u0.w[0][17] ),
    .Z(_17107_));
 CLKBUF_X1 _33940_ (.A(net49),
    .Z(_01309_));
 CLKBUF_X1 _33941_ (.A(_01098_),
    .Z(_00499_));
 CLKBUF_X2 _33942_ (.A(\u0.w[1][18] ),
    .Z(_17140_));
 CLKBUF_X2 _33943_ (.A(\u0.w[0][18] ),
    .Z(_17108_));
 CLKBUF_X1 _33944_ (.A(net48),
    .Z(_01310_));
 CLKBUF_X1 _33945_ (.A(_01099_),
    .Z(_00500_));
 CLKBUF_X2 _33946_ (.A(\u0.w[1][19] ),
    .Z(_17141_));
 CLKBUF_X2 _33947_ (.A(\u0.w[0][19] ),
    .Z(_17109_));
 CLKBUF_X1 _33948_ (.A(net47),
    .Z(_01311_));
 CLKBUF_X1 _33949_ (.A(_01100_),
    .Z(_00501_));
 CLKBUF_X2 _33950_ (.A(\u0.w[1][20] ),
    .Z(_17143_));
 BUF_X1 _33951_ (.A(\u0.w[0][20] ),
    .Z(_17111_));
 CLKBUF_X1 _33952_ (.A(net46),
    .Z(_01312_));
 CLKBUF_X1 _33953_ (.A(_01102_),
    .Z(_00503_));
 CLKBUF_X1 _33954_ (.A(\u0.w[1][21] ),
    .Z(_17144_));
 CLKBUF_X1 _33955_ (.A(\u0.w[0][21] ),
    .Z(_17112_));
 CLKBUF_X1 _33956_ (.A(net45),
    .Z(_01313_));
 CLKBUF_X1 _33957_ (.A(_01103_),
    .Z(_00504_));
 CLKBUF_X1 _33958_ (.A(\u0.w[1][22] ),
    .Z(_17145_));
 CLKBUF_X1 _33959_ (.A(\u0.w[0][22] ),
    .Z(_17113_));
 CLKBUF_X1 _33960_ (.A(net44),
    .Z(_01314_));
 CLKBUF_X1 _33961_ (.A(_01104_),
    .Z(_00505_));
 CLKBUF_X2 _33962_ (.A(\u0.w[1][23] ),
    .Z(_17146_));
 BUF_X1 _33963_ (.A(\u0.w[0][23] ),
    .Z(_17114_));
 CLKBUF_X1 _33964_ (.A(net43),
    .Z(_01315_));
 CLKBUF_X1 _33965_ (.A(_01105_),
    .Z(_00506_));
 CLKBUF_X1 _33966_ (.A(\u0.w[0][24] ),
    .Z(_17115_));
 CLKBUF_X1 _33967_ (.A(\u0.w[1][24] ),
    .Z(_17147_));
 CLKBUF_X1 _33968_ (.A(net42),
    .Z(_01316_));
 CLKBUF_X1 _33969_ (.A(_01106_),
    .Z(_00507_));
 CLKBUF_X1 _33970_ (.A(\u0.w[0][25] ),
    .Z(_17116_));
 CLKBUF_X1 _33971_ (.A(\u0.w[1][25] ),
    .Z(_17148_));
 CLKBUF_X1 _33972_ (.A(net41),
    .Z(_01317_));
 CLKBUF_X1 _33973_ (.A(_01107_),
    .Z(_00508_));
 CLKBUF_X1 _33974_ (.A(\u0.w[0][26] ),
    .Z(_17117_));
 BUF_X1 _33975_ (.A(\u0.w[1][26] ),
    .Z(_17149_));
 CLKBUF_X1 _33976_ (.A(net40),
    .Z(_01319_));
 CLKBUF_X1 _33977_ (.A(_01108_),
    .Z(_00509_));
 BUF_X1 _33978_ (.A(\u0.w[0][27] ),
    .Z(_17118_));
 BUF_X1 _33979_ (.A(\u0.w[1][27] ),
    .Z(_17150_));
 CLKBUF_X1 _33980_ (.A(net39),
    .Z(_01320_));
 CLKBUF_X1 _33981_ (.A(_01109_),
    .Z(_00510_));
 BUF_X1 _33982_ (.A(\u0.w[0][28] ),
    .Z(_17119_));
 CLKBUF_X2 _33983_ (.A(\u0.w[1][28] ),
    .Z(_17151_));
 CLKBUF_X1 _33984_ (.A(net38),
    .Z(_01321_));
 CLKBUF_X1 _33985_ (.A(_01110_),
    .Z(_00511_));
 CLKBUF_X1 _33986_ (.A(\u0.w[0][29] ),
    .Z(_17120_));
 CLKBUF_X1 _33987_ (.A(\u0.w[1][29] ),
    .Z(_17152_));
 CLKBUF_X1 _33988_ (.A(net37),
    .Z(_01322_));
 CLKBUF_X1 _33989_ (.A(_01111_),
    .Z(_00512_));
 CLKBUF_X1 _33990_ (.A(\u0.w[0][30] ),
    .Z(_17122_));
 CLKBUF_X1 _33991_ (.A(\u0.w[1][30] ),
    .Z(_17154_));
 CLKBUF_X1 _33992_ (.A(net36),
    .Z(_01323_));
 CLKBUF_X1 _33993_ (.A(_01113_),
    .Z(_00514_));
 BUF_X1 _33994_ (.A(\u0.w[0][31] ),
    .Z(_17123_));
 CLKBUF_X2 _33995_ (.A(\u0.w[1][31] ),
    .Z(_17155_));
 CLKBUF_X1 _33996_ (.A(net35),
    .Z(_01324_));
 CLKBUF_X1 _33997_ (.A(_01114_),
    .Z(_00515_));
 CLKBUF_X1 _33998_ (.A(_00430_),
    .Z(_01029_));
 CLKBUF_X1 _33999_ (.A(\u0.w[2][16] ),
    .Z(_17170_));
 CLKBUF_X1 _34000_ (.A(\text_in_r[48] ),
    .Z(_17005_));
 CLKBUF_X1 _34001_ (.A(_00652_),
    .Z(_00053_));
 CLKBUF_X1 _34002_ (.A(_00431_),
    .Z(_01030_));
 CLKBUF_X1 _34003_ (.A(\u0.w[2][17] ),
    .Z(_17171_));
 CLKBUF_X1 _34004_ (.A(\text_in_r[49] ),
    .Z(_17006_));
 CLKBUF_X1 _34005_ (.A(_00653_),
    .Z(_00054_));
 BUF_X1 _34006_ (.A(\u0.w[2][18] ),
    .Z(_17172_));
 CLKBUF_X1 _34007_ (.A(\text_in_r[50] ),
    .Z(_17008_));
 CLKBUF_X1 _34008_ (.A(_00654_),
    .Z(_00055_));
 CLKBUF_X2 _34009_ (.A(\u0.w[2][19] ),
    .Z(_17173_));
 CLKBUF_X1 _34010_ (.A(\text_in_r[51] ),
    .Z(_17009_));
 CLKBUF_X1 _34011_ (.A(_00655_),
    .Z(_00056_));
 BUF_X1 _34012_ (.A(\u0.w[2][20] ),
    .Z(_17175_));
 CLKBUF_X1 _34013_ (.A(\text_in_r[52] ),
    .Z(_17010_));
 CLKBUF_X1 _34014_ (.A(_00656_),
    .Z(_00057_));
 CLKBUF_X1 _34015_ (.A(_00432_),
    .Z(_01031_));
 CLKBUF_X1 _34016_ (.A(\u0.w[2][21] ),
    .Z(_17176_));
 CLKBUF_X1 _34017_ (.A(\text_in_r[53] ),
    .Z(_17011_));
 CLKBUF_X1 _34018_ (.A(_00657_),
    .Z(_00058_));
 CLKBUF_X1 _34019_ (.A(_00433_),
    .Z(_01032_));
 CLKBUF_X1 _34020_ (.A(\u0.w[2][22] ),
    .Z(_17177_));
 CLKBUF_X1 _34021_ (.A(\text_in_r[54] ),
    .Z(_17012_));
 CLKBUF_X1 _34022_ (.A(_00658_),
    .Z(_00059_));
 BUF_X1 _34023_ (.A(\u0.w[2][23] ),
    .Z(_17178_));
 CLKBUF_X1 _34024_ (.A(\text_in_r[55] ),
    .Z(_17013_));
 CLKBUF_X1 _34025_ (.A(_00659_),
    .Z(_00060_));
 CLKBUF_X1 _34026_ (.A(net98),
    .Z(_01255_));
 CLKBUF_X1 _34027_ (.A(_01122_),
    .Z(_00523_));
 CLKBUF_X1 _34028_ (.A(net97),
    .Z(_01256_));
 CLKBUF_X1 _34029_ (.A(_01133_),
    .Z(_00534_));
 CLKBUF_X1 _34030_ (.A(net96),
    .Z(_01257_));
 CLKBUF_X1 _34031_ (.A(_01144_),
    .Z(_00545_));
 CLKBUF_X1 _34032_ (.A(net95),
    .Z(_01258_));
 CLKBUF_X1 _34033_ (.A(_01147_),
    .Z(_00548_));
 CLKBUF_X1 _34034_ (.A(net94),
    .Z(_01259_));
 CLKBUF_X1 _34035_ (.A(_01148_),
    .Z(_00549_));
 CLKBUF_X1 _34036_ (.A(net93),
    .Z(_01260_));
 CLKBUF_X1 _34037_ (.A(_01149_),
    .Z(_00550_));
 CLKBUF_X1 _34038_ (.A(net92),
    .Z(_01261_));
 CLKBUF_X1 _34039_ (.A(_01150_),
    .Z(_00551_));
 CLKBUF_X1 _34040_ (.A(net91),
    .Z(_01262_));
 CLKBUF_X1 _34041_ (.A(_01151_),
    .Z(_00552_));
 CLKBUF_X1 _34042_ (.A(net90),
    .Z(_01264_));
 CLKBUF_X1 _34043_ (.A(_01152_),
    .Z(_00553_));
 CLKBUF_X1 _34044_ (.A(net89),
    .Z(_01265_));
 CLKBUF_X1 _34045_ (.A(_01153_),
    .Z(_00554_));
 CLKBUF_X1 _34046_ (.A(net88),
    .Z(_01266_));
 CLKBUF_X1 _34047_ (.A(_01123_),
    .Z(_00524_));
 CLKBUF_X1 _34048_ (.A(net87),
    .Z(_01267_));
 CLKBUF_X1 _34049_ (.A(_01124_),
    .Z(_00525_));
 CLKBUF_X1 _34050_ (.A(net86),
    .Z(_01268_));
 CLKBUF_X1 _34051_ (.A(_01125_),
    .Z(_00526_));
 CLKBUF_X1 _34052_ (.A(net85),
    .Z(_01269_));
 CLKBUF_X1 _34053_ (.A(_01126_),
    .Z(_00527_));
 CLKBUF_X1 _34054_ (.A(net84),
    .Z(_01270_));
 CLKBUF_X1 _34055_ (.A(_01127_),
    .Z(_00528_));
 CLKBUF_X1 _34056_ (.A(net83),
    .Z(_01271_));
 CLKBUF_X1 _34057_ (.A(_01128_),
    .Z(_00529_));
 CLKBUF_X1 _34058_ (.A(net82),
    .Z(_01272_));
 CLKBUF_X1 _34059_ (.A(_01129_),
    .Z(_00530_));
 CLKBUF_X1 _34060_ (.A(net81),
    .Z(_01273_));
 CLKBUF_X1 _34061_ (.A(_01130_),
    .Z(_00531_));
 CLKBUF_X1 _34062_ (.A(net80),
    .Z(_01275_));
 CLKBUF_X1 _34063_ (.A(_01131_),
    .Z(_00532_));
 CLKBUF_X1 _34064_ (.A(net79),
    .Z(_01276_));
 CLKBUF_X1 _34065_ (.A(_01132_),
    .Z(_00533_));
 CLKBUF_X1 _34066_ (.A(net78),
    .Z(_01277_));
 CLKBUF_X1 _34067_ (.A(_01134_),
    .Z(_00535_));
 CLKBUF_X1 _34068_ (.A(net77),
    .Z(_01278_));
 CLKBUF_X1 _34069_ (.A(_01135_),
    .Z(_00536_));
 CLKBUF_X1 _34070_ (.A(net76),
    .Z(_01279_));
 CLKBUF_X1 _34071_ (.A(_01136_),
    .Z(_00537_));
 CLKBUF_X1 _34072_ (.A(net75),
    .Z(_01280_));
 CLKBUF_X1 _34073_ (.A(_01137_),
    .Z(_00538_));
 CLKBUF_X1 _34074_ (.A(\u0.w[2][24] ),
    .Z(_17179_));
 CLKBUF_X1 _34075_ (.A(net74),
    .Z(_01281_));
 CLKBUF_X1 _34076_ (.A(_01138_),
    .Z(_00539_));
 CLKBUF_X1 _34077_ (.A(\u0.w[2][25] ),
    .Z(_17180_));
 CLKBUF_X1 _34078_ (.A(net73),
    .Z(_01282_));
 CLKBUF_X1 _34079_ (.A(_01139_),
    .Z(_00540_));
 CLKBUF_X2 _34080_ (.A(\u0.w[2][26] ),
    .Z(_17181_));
 CLKBUF_X1 _34081_ (.A(net72),
    .Z(_01283_));
 CLKBUF_X1 _34082_ (.A(_01140_),
    .Z(_00541_));
 CLKBUF_X2 _34083_ (.A(\u0.w[2][27] ),
    .Z(_17182_));
 CLKBUF_X1 _34084_ (.A(net71),
    .Z(_01284_));
 CLKBUF_X1 _34085_ (.A(_01141_),
    .Z(_00542_));
 CLKBUF_X2 _34086_ (.A(\u0.w[2][28] ),
    .Z(_17183_));
 CLKBUF_X1 _34087_ (.A(net70),
    .Z(_01286_));
 CLKBUF_X1 _34088_ (.A(_01142_),
    .Z(_00543_));
 CLKBUF_X1 _34089_ (.A(\u0.w[2][29] ),
    .Z(_17184_));
 CLKBUF_X1 _34090_ (.A(net69),
    .Z(_01287_));
 CLKBUF_X1 _34091_ (.A(_01143_),
    .Z(_00544_));
 CLKBUF_X1 _34092_ (.A(\u0.w[2][30] ),
    .Z(_17186_));
 CLKBUF_X1 _34093_ (.A(net68),
    .Z(_01288_));
 CLKBUF_X1 _34094_ (.A(_01145_),
    .Z(_00546_));
 BUF_X1 _34095_ (.A(\u0.w[2][31] ),
    .Z(_17187_));
 CLKBUF_X1 _34096_ (.A(net67),
    .Z(_01289_));
 CLKBUF_X1 _34097_ (.A(_01146_),
    .Z(_00547_));
 CLKBUF_X1 _34098_ (.A(_00434_),
    .Z(_01033_));
 CLKBUF_X1 _34099_ (.A(\text_in_r[56] ),
    .Z(_17014_));
 CLKBUF_X1 _34100_ (.A(_00620_),
    .Z(_00021_));
 CLKBUF_X1 _34101_ (.A(_00435_),
    .Z(_01034_));
 CLKBUF_X1 _34102_ (.A(\text_in_r[57] ),
    .Z(_17015_));
 CLKBUF_X1 _34103_ (.A(_00621_),
    .Z(_00022_));
 CLKBUF_X1 _34104_ (.A(\text_in_r[58] ),
    .Z(_17016_));
 CLKBUF_X1 _34105_ (.A(_00622_),
    .Z(_00023_));
 CLKBUF_X1 _34106_ (.A(\text_in_r[59] ),
    .Z(_17017_));
 CLKBUF_X1 _34107_ (.A(_00623_),
    .Z(_00024_));
 CLKBUF_X1 _34108_ (.A(\text_in_r[60] ),
    .Z(_17019_));
 CLKBUF_X1 _34109_ (.A(_00624_),
    .Z(_00025_));
 CLKBUF_X1 _34110_ (.A(_00436_),
    .Z(_01035_));
 CLKBUF_X1 _34111_ (.A(\text_in_r[61] ),
    .Z(_17020_));
 CLKBUF_X1 _34112_ (.A(_00625_),
    .Z(_00026_));
 CLKBUF_X1 _34113_ (.A(_00437_),
    .Z(_01036_));
 CLKBUF_X1 _34114_ (.A(\text_in_r[62] ),
    .Z(_17021_));
 CLKBUF_X1 _34115_ (.A(_00626_),
    .Z(_00027_));
 CLKBUF_X1 _34116_ (.A(\text_in_r[63] ),
    .Z(_17022_));
 CLKBUF_X1 _34117_ (.A(_00627_),
    .Z(_00028_));
 CLKBUF_X1 _34118_ (.A(net130),
    .Z(_01202_));
 CLKBUF_X1 _34119_ (.A(_01154_),
    .Z(_00555_));
 CLKBUF_X1 _34120_ (.A(net129),
    .Z(_01241_));
 CLKBUF_X1 _34121_ (.A(_01165_),
    .Z(_00566_));
 CLKBUF_X1 _34122_ (.A(\sa01[5] ),
    .Z(_16692_));
 CLKBUF_X1 _34123_ (.A(\sa01[4] ),
    .Z(_16691_));
 CLKBUF_X1 _34124_ (.A(\sa01[7] ),
    .Z(_16694_));
 BUF_X1 _34125_ (.A(\sa01[6] ),
    .Z(_16693_));
 CLKBUF_X2 _34126_ (.A(\sa01[1] ),
    .Z(_16688_));
 CLKBUF_X2 _34127_ (.A(\sa01[0] ),
    .Z(_16687_));
 CLKBUF_X2 _34128_ (.A(\sa01[2] ),
    .Z(_16689_));
 CLKBUF_X2 _34129_ (.A(\sa01[3] ),
    .Z(_16690_));
 CLKBUF_X1 _34130_ (.A(\sa12[5] ),
    .Z(_16732_));
 BUF_X1 _34131_ (.A(\sa12[4] ),
    .Z(_16731_));
 CLKBUF_X1 _34132_ (.A(\sa12[7] ),
    .Z(_16734_));
 CLKBUF_X1 _34133_ (.A(\sa12[6] ),
    .Z(_16733_));
 CLKBUF_X2 _34134_ (.A(\sa12[1] ),
    .Z(_16728_));
 BUF_X1 _34135_ (.A(\sa12[0] ),
    .Z(_16727_));
 BUF_X1 _34136_ (.A(\sa12[2] ),
    .Z(_16729_));
 CLKBUF_X2 _34137_ (.A(\sa12[3] ),
    .Z(_16730_));
 CLKBUF_X1 _34138_ (.A(\sa23[5] ),
    .Z(_16772_));
 CLKBUF_X1 _34139_ (.A(\sa23[4] ),
    .Z(_16771_));
 CLKBUF_X1 _34140_ (.A(\sa23[7] ),
    .Z(_16774_));
 CLKBUF_X1 _34141_ (.A(\sa23[6] ),
    .Z(_16773_));
 BUF_X1 _34142_ (.A(\sa23[1] ),
    .Z(_16768_));
 CLKBUF_X1 _34143_ (.A(\sa23[0] ),
    .Z(_16767_));
 CLKBUF_X2 _34144_ (.A(\sa23[2] ),
    .Z(_16769_));
 CLKBUF_X2 _34145_ (.A(\sa23[3] ),
    .Z(_16770_));
 CLKBUF_X1 _34146_ (.A(\sa30[0] ),
    .Z(_16775_));
 BUF_X1 _34147_ (.A(\sa30[1] ),
    .Z(_16776_));
 BUF_X1 _34148_ (.A(\sa30[2] ),
    .Z(_16777_));
 CLKBUF_X2 _34149_ (.A(\sa30[3] ),
    .Z(_16778_));
 BUF_X1 _34150_ (.A(\sa30[5] ),
    .Z(_16780_));
 BUF_X1 _34151_ (.A(\sa30[4] ),
    .Z(_16779_));
 CLKBUF_X1 _34152_ (.A(\sa30[7] ),
    .Z(_16782_));
 CLKBUF_X1 _34153_ (.A(\sa30[6] ),
    .Z(_16781_));
 CLKBUF_X1 _34154_ (.A(\text_in_r[64] ),
    .Z(_17023_));
 CLKBUF_X1 _34155_ (.A(_00708_),
    .Z(_00109_));
 CLKBUF_X1 _34156_ (.A(net128),
    .Z(_01252_));
 CLKBUF_X1 _34157_ (.A(_01176_),
    .Z(_00577_));
 CLKBUF_X1 _34158_ (.A(net127),
    .Z(_01263_));
 CLKBUF_X1 _34159_ (.A(_01179_),
    .Z(_00580_));
 CLKBUF_X1 _34160_ (.A(net126),
    .Z(_01274_));
 CLKBUF_X1 _34161_ (.A(_01180_),
    .Z(_00581_));
 CLKBUF_X1 _34162_ (.A(net125),
    .Z(_01285_));
 CLKBUF_X1 _34163_ (.A(_01181_),
    .Z(_00582_));
 CLKBUF_X1 _34164_ (.A(net124),
    .Z(_01296_));
 CLKBUF_X1 _34165_ (.A(_01182_),
    .Z(_00583_));
 CLKBUF_X1 _34166_ (.A(net123),
    .Z(_01307_));
 CLKBUF_X1 _34167_ (.A(_01183_),
    .Z(_00584_));
 CLKBUF_X1 _34168_ (.A(net122),
    .Z(_01318_));
 CLKBUF_X1 _34169_ (.A(_01184_),
    .Z(_00585_));
 CLKBUF_X1 _34170_ (.A(net121),
    .Z(_01329_));
 CLKBUF_X1 _34171_ (.A(_01185_),
    .Z(_00586_));
 CLKBUF_X1 _34172_ (.A(net120),
    .Z(_01213_));
 CLKBUF_X1 _34173_ (.A(_01155_),
    .Z(_00556_));
 CLKBUF_X1 _34174_ (.A(net119),
    .Z(_01224_));
 CLKBUF_X1 _34175_ (.A(_01156_),
    .Z(_00557_));
 CLKBUF_X1 _34176_ (.A(\text_in_r[65] ),
    .Z(_17024_));
 CLKBUF_X1 _34177_ (.A(_00709_),
    .Z(_00110_));
 CLKBUF_X1 _34178_ (.A(net118),
    .Z(_01233_));
 CLKBUF_X1 _34179_ (.A(_01157_),
    .Z(_00558_));
 CLKBUF_X1 _34180_ (.A(net117),
    .Z(_01234_));
 CLKBUF_X1 _34181_ (.A(_01158_),
    .Z(_00559_));
 CLKBUF_X1 _34182_ (.A(net116),
    .Z(_01235_));
 CLKBUF_X1 _34183_ (.A(_01159_),
    .Z(_00560_));
 CLKBUF_X1 _34184_ (.A(net115),
    .Z(_01236_));
 CLKBUF_X1 _34185_ (.A(_01160_),
    .Z(_00561_));
 CLKBUF_X1 _34186_ (.A(net114),
    .Z(_01237_));
 CLKBUF_X1 _34187_ (.A(_01161_),
    .Z(_00562_));
 CLKBUF_X1 _34188_ (.A(net113),
    .Z(_01238_));
 CLKBUF_X1 _34189_ (.A(_01162_),
    .Z(_00563_));
 CLKBUF_X1 _34190_ (.A(net112),
    .Z(_01239_));
 CLKBUF_X1 _34191_ (.A(_01163_),
    .Z(_00564_));
 CLKBUF_X1 _34192_ (.A(net111),
    .Z(_01240_));
 CLKBUF_X1 _34193_ (.A(_01164_),
    .Z(_00565_));
 CLKBUF_X1 _34194_ (.A(net110),
    .Z(_01242_));
 CLKBUF_X1 _34195_ (.A(_01166_),
    .Z(_00567_));
 CLKBUF_X1 _34196_ (.A(net109),
    .Z(_01243_));
 CLKBUF_X1 _34197_ (.A(_01167_),
    .Z(_00568_));
 CLKBUF_X1 _34198_ (.A(\text_in_r[66] ),
    .Z(_17025_));
 CLKBUF_X1 _34199_ (.A(_00710_),
    .Z(_00111_));
 CLKBUF_X1 _34200_ (.A(net108),
    .Z(_01244_));
 CLKBUF_X1 _34201_ (.A(_01168_),
    .Z(_00569_));
 CLKBUF_X1 _34202_ (.A(net107),
    .Z(_01245_));
 CLKBUF_X1 _34203_ (.A(_01169_),
    .Z(_00570_));
 CLKBUF_X1 _34204_ (.A(net106),
    .Z(_01246_));
 CLKBUF_X1 _34205_ (.A(_01170_),
    .Z(_00571_));
 CLKBUF_X1 _34206_ (.A(net105),
    .Z(_01247_));
 CLKBUF_X1 _34207_ (.A(_01171_),
    .Z(_00572_));
 CLKBUF_X1 _34208_ (.A(net104),
    .Z(_01248_));
 CLKBUF_X1 _34209_ (.A(_01172_),
    .Z(_00573_));
 CLKBUF_X1 _34210_ (.A(net103),
    .Z(_01249_));
 CLKBUF_X1 _34211_ (.A(_01173_),
    .Z(_00574_));
 CLKBUF_X1 _34212_ (.A(net102),
    .Z(_01250_));
 CLKBUF_X1 _34213_ (.A(_01174_),
    .Z(_00575_));
 CLKBUF_X1 _34214_ (.A(net101),
    .Z(_01251_));
 CLKBUF_X1 _34215_ (.A(_01175_),
    .Z(_00576_));
 CLKBUF_X1 _34216_ (.A(net100),
    .Z(_01253_));
 CLKBUF_X1 _34217_ (.A(_01177_),
    .Z(_00578_));
 CLKBUF_X1 _34218_ (.A(net99),
    .Z(_01254_));
 CLKBUF_X1 _34219_ (.A(_01178_),
    .Z(_00579_));
 CLKBUF_X1 _34220_ (.A(\text_in_r[67] ),
    .Z(_17026_));
 CLKBUF_X1 _34221_ (.A(_00711_),
    .Z(_00112_));
 CLKBUF_X1 _34222_ (.A(\text_in_r[68] ),
    .Z(_17027_));
 CLKBUF_X1 _34223_ (.A(_00712_),
    .Z(_00113_));
 CLKBUF_X1 _34224_ (.A(\text_in_r[69] ),
    .Z(_17028_));
 CLKBUF_X1 _34225_ (.A(_00713_),
    .Z(_00114_));
 CLKBUF_X1 _34226_ (.A(\text_in_r[70] ),
    .Z(_17030_));
 CLKBUF_X1 _34227_ (.A(_00714_),
    .Z(_00115_));
 CLKBUF_X1 _34228_ (.A(\text_in_r[71] ),
    .Z(_17031_));
 CLKBUF_X1 _34229_ (.A(_00715_),
    .Z(_00116_));
 CLKBUF_X1 _34230_ (.A(_00438_),
    .Z(_01037_));
 CLKBUF_X1 _34231_ (.A(\text_in_r[72] ),
    .Z(_17032_));
 CLKBUF_X1 _34232_ (.A(_00676_),
    .Z(_00077_));
 CLKBUF_X1 _34233_ (.A(\text_in_r[73] ),
    .Z(_17033_));
 CLKBUF_X1 _34234_ (.A(_00677_),
    .Z(_00078_));
 CLKBUF_X1 _34235_ (.A(\text_in_r[74] ),
    .Z(_17034_));
 CLKBUF_X1 _34236_ (.A(_00678_),
    .Z(_00079_));
 CLKBUF_X1 _34237_ (.A(\text_in_r[75] ),
    .Z(_17035_));
 CLKBUF_X1 _34238_ (.A(_00679_),
    .Z(_00080_));
 CLKBUF_X1 _34239_ (.A(\text_in_r[76] ),
    .Z(_17036_));
 CLKBUF_X1 _34240_ (.A(_00680_),
    .Z(_00081_));
 CLKBUF_X1 _34241_ (.A(\text_in_r[77] ),
    .Z(_17037_));
 CLKBUF_X1 _34242_ (.A(_00681_),
    .Z(_00082_));
 CLKBUF_X1 _34243_ (.A(\text_in_r[78] ),
    .Z(_17038_));
 CLKBUF_X1 _34244_ (.A(_00682_),
    .Z(_00083_));
 CLKBUF_X1 _34245_ (.A(\text_in_r[79] ),
    .Z(_17039_));
 CLKBUF_X1 _34246_ (.A(_00683_),
    .Z(_00084_));
 CLKBUF_X1 _34247_ (.A(_00439_),
    .Z(_01038_));
 CLKBUF_X1 _34248_ (.A(\text_in_r[80] ),
    .Z(_17041_));
 CLKBUF_X1 _34249_ (.A(_00644_),
    .Z(_00045_));
 CLKBUF_X1 _34250_ (.A(_00440_),
    .Z(_01039_));
 CLKBUF_X1 _34251_ (.A(\text_in_r[81] ),
    .Z(_17042_));
 CLKBUF_X1 _34252_ (.A(_00645_),
    .Z(_00046_));
 CLKBUF_X1 _34253_ (.A(\text_in_r[82] ),
    .Z(_17043_));
 CLKBUF_X1 _34254_ (.A(_00646_),
    .Z(_00047_));
 CLKBUF_X1 _34255_ (.A(\text_in_r[83] ),
    .Z(_17044_));
 CLKBUF_X1 _34256_ (.A(_00647_),
    .Z(_00048_));
 CLKBUF_X1 _34257_ (.A(\text_in_r[84] ),
    .Z(_17045_));
 CLKBUF_X1 _34258_ (.A(_00648_),
    .Z(_00049_));
 CLKBUF_X1 _34259_ (.A(_00441_),
    .Z(_01040_));
 CLKBUF_X1 _34260_ (.A(\text_in_r[85] ),
    .Z(_17046_));
 CLKBUF_X1 _34261_ (.A(_00649_),
    .Z(_00050_));
 CLKBUF_X1 _34262_ (.A(_00442_),
    .Z(_01041_));
 CLKBUF_X1 _34263_ (.A(\text_in_r[86] ),
    .Z(_17047_));
 CLKBUF_X1 _34264_ (.A(_00650_),
    .Z(_00051_));
 CLKBUF_X1 _34265_ (.A(\text_in_r[87] ),
    .Z(_17048_));
 CLKBUF_X1 _34266_ (.A(_00651_),
    .Z(_00052_));
 CLKBUF_X1 _34267_ (.A(_00443_),
    .Z(_01042_));
 CLKBUF_X1 _34268_ (.A(\text_in_r[88] ),
    .Z(_17049_));
 CLKBUF_X1 _34269_ (.A(_00612_),
    .Z(_00013_));
 CLKBUF_X1 _34270_ (.A(_00444_),
    .Z(_01043_));
 CLKBUF_X1 _34271_ (.A(\text_in_r[89] ),
    .Z(_17050_));
 CLKBUF_X1 _34272_ (.A(_00613_),
    .Z(_00014_));
 CLKBUF_X1 _34273_ (.A(\text_in_r[90] ),
    .Z(_17052_));
 CLKBUF_X1 _34274_ (.A(_00614_),
    .Z(_00015_));
 CLKBUF_X1 _34275_ (.A(\text_in_r[91] ),
    .Z(_17053_));
 CLKBUF_X1 _34276_ (.A(_00615_),
    .Z(_00016_));
 CLKBUF_X1 _34277_ (.A(\text_in_r[92] ),
    .Z(_17054_));
 CLKBUF_X1 _34278_ (.A(_00616_),
    .Z(_00017_));
 CLKBUF_X1 _34279_ (.A(_00445_),
    .Z(_01044_));
 CLKBUF_X1 _34280_ (.A(\text_in_r[93] ),
    .Z(_17055_));
 CLKBUF_X1 _34281_ (.A(_00617_),
    .Z(_00018_));
 CLKBUF_X1 _34282_ (.A(net1),
    .Z(_16678_));
 CLKBUF_X1 _34283_ (.A(\dcnt[2] ),
    .Z(_01200_));
 CLKBUF_X1 _34284_ (.A(\dcnt[3] ),
    .Z(_01201_));
 CLKBUF_X1 _34285_ (.A(\dcnt[0] ),
    .Z(_01198_));
 CLKBUF_X1 _34286_ (.A(\dcnt[1] ),
    .Z(_01199_));
 CLKBUF_X1 _34287_ (.A(_00599_),
    .Z(_00000_));
 CLKBUF_X1 _34288_ (.A(_00446_),
    .Z(_01045_));
 CLKBUF_X1 _34289_ (.A(_00600_),
    .Z(_00001_));
 CLKBUF_X1 _34290_ (.A(_00447_),
    .Z(_01046_));
 CLKBUF_X1 _34291_ (.A(_00601_),
    .Z(_00002_));
 CLKBUF_X1 _34292_ (.A(_00448_),
    .Z(_01047_));
 CLKBUF_X1 _34293_ (.A(_00602_),
    .Z(_00003_));
 CLKBUF_X1 _34294_ (.A(_00449_),
    .Z(_01048_));
 CLKBUF_X1 _34295_ (.A(\text_in_r[94] ),
    .Z(_17056_));
 CLKBUF_X1 _34296_ (.A(_00618_),
    .Z(_00019_));
 CLKBUF_X1 _34297_ (.A(net258),
    .Z(_16807_));
 CLKBUF_X1 _34298_ (.A(_00732_),
    .Z(_00133_));
 CLKBUF_X1 _34299_ (.A(net257),
    .Z(_16846_));
 CLKBUF_X1 _34300_ (.A(_00771_),
    .Z(_00172_));
 CLKBUF_X1 _34301_ (.A(net256),
    .Z(_16857_));
 CLKBUF_X1 _34302_ (.A(_00782_),
    .Z(_00183_));
 CLKBUF_X1 _34303_ (.A(net255),
    .Z(_16868_));
 CLKBUF_X1 _34304_ (.A(_00793_),
    .Z(_00194_));
 CLKBUF_X1 _34305_ (.A(net254),
    .Z(_16879_));
 CLKBUF_X1 _34306_ (.A(_00804_),
    .Z(_00205_));
 CLKBUF_X1 _34307_ (.A(net253),
    .Z(_16890_));
 CLKBUF_X1 _34308_ (.A(_00815_),
    .Z(_00216_));
 CLKBUF_X1 _34309_ (.A(\text_in_r[95] ),
    .Z(_17057_));
 CLKBUF_X1 _34310_ (.A(_00619_),
    .Z(_00020_));
 CLKBUF_X1 _34311_ (.A(net252),
    .Z(_16901_));
 CLKBUF_X1 _34312_ (.A(_00826_),
    .Z(_00227_));
 CLKBUF_X1 _34313_ (.A(net251),
    .Z(_16912_));
 CLKBUF_X1 _34314_ (.A(_00837_),
    .Z(_00238_));
 CLKBUF_X1 _34315_ (.A(net250),
    .Z(_16923_));
 CLKBUF_X1 _34316_ (.A(_00848_),
    .Z(_00249_));
 CLKBUF_X1 _34317_ (.A(net249),
    .Z(_16934_));
 CLKBUF_X1 _34318_ (.A(_00859_),
    .Z(_00260_));
 CLKBUF_X1 _34319_ (.A(net248),
    .Z(_16818_));
 CLKBUF_X1 _34320_ (.A(_00743_),
    .Z(_00144_));
 CLKBUF_X1 _34321_ (.A(net247),
    .Z(_16829_));
 CLKBUF_X1 _34322_ (.A(_00754_),
    .Z(_00155_));
 CLKBUF_X1 _34323_ (.A(net246),
    .Z(_16838_));
 CLKBUF_X1 _34324_ (.A(_00763_),
    .Z(_00164_));
 CLKBUF_X1 _34325_ (.A(net245),
    .Z(_16839_));
 CLKBUF_X1 _34326_ (.A(_00764_),
    .Z(_00165_));
 CLKBUF_X1 _34327_ (.A(net244),
    .Z(_16840_));
 CLKBUF_X1 _34328_ (.A(_00765_),
    .Z(_00166_));
 CLKBUF_X1 _34329_ (.A(net243),
    .Z(_16841_));
 CLKBUF_X1 _34330_ (.A(_00766_),
    .Z(_00167_));
 CLKBUF_X1 _34331_ (.A(net242),
    .Z(_16842_));
 CLKBUF_X1 _34332_ (.A(_00767_),
    .Z(_00168_));
 CLKBUF_X1 _34333_ (.A(net241),
    .Z(_16843_));
 CLKBUF_X1 _34334_ (.A(_00768_),
    .Z(_00169_));
 CLKBUF_X1 _34335_ (.A(net240),
    .Z(_16844_));
 CLKBUF_X1 _34336_ (.A(_00769_),
    .Z(_00170_));
 CLKBUF_X1 _34337_ (.A(net239),
    .Z(_16845_));
 CLKBUF_X1 _34338_ (.A(_00770_),
    .Z(_00171_));
 CLKBUF_X1 _34339_ (.A(net238),
    .Z(_16847_));
 CLKBUF_X1 _34340_ (.A(_00772_),
    .Z(_00173_));
 CLKBUF_X1 _34341_ (.A(net237),
    .Z(_16848_));
 CLKBUF_X1 _34342_ (.A(_00773_),
    .Z(_00174_));
 CLKBUF_X1 _34343_ (.A(net236),
    .Z(_16849_));
 CLKBUF_X1 _34344_ (.A(_00774_),
    .Z(_00175_));
 CLKBUF_X1 _34345_ (.A(net235),
    .Z(_16850_));
 CLKBUF_X1 _34346_ (.A(_00775_),
    .Z(_00176_));
 CLKBUF_X1 _34347_ (.A(net234),
    .Z(_16851_));
 CLKBUF_X1 _34348_ (.A(_00776_),
    .Z(_00177_));
 CLKBUF_X1 _34349_ (.A(net233),
    .Z(_16852_));
 CLKBUF_X1 _34350_ (.A(_00777_),
    .Z(_00178_));
 CLKBUF_X1 _34351_ (.A(net232),
    .Z(_16853_));
 CLKBUF_X1 _34352_ (.A(_00778_),
    .Z(_00179_));
 CLKBUF_X1 _34353_ (.A(net231),
    .Z(_16854_));
 CLKBUF_X1 _34354_ (.A(_00779_),
    .Z(_00180_));
 CLKBUF_X1 _34355_ (.A(net230),
    .Z(_16855_));
 CLKBUF_X1 _34356_ (.A(_00780_),
    .Z(_00181_));
 CLKBUF_X1 _34357_ (.A(net229),
    .Z(_16856_));
 CLKBUF_X1 _34358_ (.A(_00781_),
    .Z(_00182_));
 CLKBUF_X1 _34359_ (.A(net228),
    .Z(_16858_));
 CLKBUF_X1 _34360_ (.A(_00783_),
    .Z(_00184_));
 CLKBUF_X1 _34361_ (.A(net227),
    .Z(_16859_));
 CLKBUF_X1 _34362_ (.A(_00784_),
    .Z(_00185_));
 CLKBUF_X1 _34363_ (.A(net226),
    .Z(_16860_));
 CLKBUF_X1 _34364_ (.A(_00785_),
    .Z(_00186_));
 CLKBUF_X1 _34365_ (.A(net225),
    .Z(_16861_));
 CLKBUF_X1 _34366_ (.A(_00786_),
    .Z(_00187_));
 CLKBUF_X1 _34367_ (.A(net224),
    .Z(_16862_));
 CLKBUF_X1 _34368_ (.A(_00787_),
    .Z(_00188_));
 CLKBUF_X1 _34369_ (.A(net223),
    .Z(_16863_));
 CLKBUF_X1 _34370_ (.A(_00788_),
    .Z(_00189_));
 CLKBUF_X1 _34371_ (.A(net222),
    .Z(_16864_));
 CLKBUF_X1 _34372_ (.A(_00789_),
    .Z(_00190_));
 CLKBUF_X1 _34373_ (.A(net221),
    .Z(_16865_));
 CLKBUF_X1 _34374_ (.A(_00790_),
    .Z(_00191_));
 CLKBUF_X1 _34375_ (.A(net220),
    .Z(_16866_));
 CLKBUF_X1 _34376_ (.A(_00791_),
    .Z(_00192_));
 CLKBUF_X1 _34377_ (.A(net219),
    .Z(_16867_));
 CLKBUF_X1 _34378_ (.A(_00792_),
    .Z(_00193_));
 CLKBUF_X1 _34379_ (.A(net218),
    .Z(_16869_));
 CLKBUF_X1 _34380_ (.A(_00794_),
    .Z(_00195_));
 CLKBUF_X1 _34381_ (.A(net217),
    .Z(_16870_));
 CLKBUF_X1 _34382_ (.A(_00795_),
    .Z(_00196_));
 CLKBUF_X1 _34383_ (.A(net216),
    .Z(_16871_));
 CLKBUF_X1 _34384_ (.A(_00796_),
    .Z(_00197_));
 CLKBUF_X1 _34385_ (.A(net215),
    .Z(_16872_));
 CLKBUF_X1 _34386_ (.A(_00797_),
    .Z(_00198_));
 CLKBUF_X1 _34387_ (.A(net214),
    .Z(_16873_));
 CLKBUF_X1 _34388_ (.A(_00798_),
    .Z(_00199_));
 CLKBUF_X1 _34389_ (.A(net213),
    .Z(_16874_));
 CLKBUF_X1 _34390_ (.A(_00799_),
    .Z(_00200_));
 CLKBUF_X1 _34391_ (.A(net212),
    .Z(_16875_));
 CLKBUF_X1 _34392_ (.A(_00800_),
    .Z(_00201_));
 CLKBUF_X1 _34393_ (.A(net211),
    .Z(_16876_));
 CLKBUF_X1 _34394_ (.A(_00801_),
    .Z(_00202_));
 CLKBUF_X1 _34395_ (.A(net210),
    .Z(_16877_));
 CLKBUF_X1 _34396_ (.A(_00802_),
    .Z(_00203_));
 CLKBUF_X1 _34397_ (.A(net209),
    .Z(_16878_));
 CLKBUF_X1 _34398_ (.A(_00803_),
    .Z(_00204_));
 CLKBUF_X1 _34399_ (.A(net208),
    .Z(_16880_));
 CLKBUF_X1 _34400_ (.A(_00805_),
    .Z(_00206_));
 CLKBUF_X1 _34401_ (.A(net207),
    .Z(_16881_));
 CLKBUF_X1 _34402_ (.A(_00806_),
    .Z(_00207_));
 CLKBUF_X1 _34403_ (.A(net206),
    .Z(_16882_));
 CLKBUF_X1 _34404_ (.A(_00807_),
    .Z(_00208_));
 CLKBUF_X1 _34405_ (.A(net205),
    .Z(_16883_));
 CLKBUF_X1 _34406_ (.A(_00808_),
    .Z(_00209_));
 CLKBUF_X1 _34407_ (.A(net204),
    .Z(_16884_));
 CLKBUF_X1 _34408_ (.A(_00809_),
    .Z(_00210_));
 CLKBUF_X1 _34409_ (.A(net203),
    .Z(_16885_));
 CLKBUF_X1 _34410_ (.A(_00810_),
    .Z(_00211_));
 CLKBUF_X1 _34411_ (.A(net202),
    .Z(_16886_));
 CLKBUF_X1 _34412_ (.A(_00811_),
    .Z(_00212_));
 CLKBUF_X1 _34413_ (.A(net201),
    .Z(_16887_));
 CLKBUF_X1 _34414_ (.A(_00812_),
    .Z(_00213_));
 CLKBUF_X1 _34415_ (.A(net200),
    .Z(_16888_));
 CLKBUF_X1 _34416_ (.A(_00813_),
    .Z(_00214_));
 CLKBUF_X1 _34417_ (.A(net199),
    .Z(_16889_));
 CLKBUF_X1 _34418_ (.A(_00814_),
    .Z(_00215_));
 CLKBUF_X1 _34419_ (.A(net198),
    .Z(_16891_));
 CLKBUF_X1 _34420_ (.A(_00816_),
    .Z(_00217_));
 CLKBUF_X1 _34421_ (.A(net197),
    .Z(_16892_));
 CLKBUF_X1 _34422_ (.A(_00817_),
    .Z(_00218_));
 CLKBUF_X1 _34423_ (.A(net196),
    .Z(_16893_));
 CLKBUF_X1 _34424_ (.A(_00818_),
    .Z(_00219_));
 CLKBUF_X1 _34425_ (.A(net195),
    .Z(_16894_));
 CLKBUF_X1 _34426_ (.A(_00819_),
    .Z(_00220_));
 CLKBUF_X1 _34427_ (.A(net194),
    .Z(_16895_));
 CLKBUF_X1 _34428_ (.A(_00820_),
    .Z(_00221_));
 CLKBUF_X1 _34429_ (.A(net193),
    .Z(_16896_));
 CLKBUF_X1 _34430_ (.A(_00821_),
    .Z(_00222_));
 CLKBUF_X1 _34431_ (.A(net192),
    .Z(_16897_));
 CLKBUF_X1 _34432_ (.A(_00822_),
    .Z(_00223_));
 CLKBUF_X1 _34433_ (.A(net191),
    .Z(_16898_));
 CLKBUF_X1 _34434_ (.A(_00823_),
    .Z(_00224_));
 CLKBUF_X1 _34435_ (.A(net190),
    .Z(_16899_));
 CLKBUF_X1 _34436_ (.A(_00824_),
    .Z(_00225_));
 CLKBUF_X1 _34437_ (.A(net189),
    .Z(_16900_));
 CLKBUF_X1 _34438_ (.A(_00825_),
    .Z(_00226_));
 CLKBUF_X1 _34439_ (.A(net188),
    .Z(_16902_));
 CLKBUF_X1 _34440_ (.A(_00827_),
    .Z(_00228_));
 CLKBUF_X1 _34441_ (.A(net187),
    .Z(_16903_));
 CLKBUF_X1 _34442_ (.A(_00828_),
    .Z(_00229_));
 CLKBUF_X1 _34443_ (.A(net186),
    .Z(_16904_));
 CLKBUF_X1 _34444_ (.A(_00829_),
    .Z(_00230_));
 CLKBUF_X1 _34445_ (.A(net185),
    .Z(_16905_));
 CLKBUF_X1 _34446_ (.A(_00830_),
    .Z(_00231_));
 CLKBUF_X1 _34447_ (.A(net184),
    .Z(_16906_));
 CLKBUF_X1 _34448_ (.A(_00831_),
    .Z(_00232_));
 CLKBUF_X1 _34449_ (.A(net183),
    .Z(_16907_));
 CLKBUF_X1 _34450_ (.A(_00832_),
    .Z(_00233_));
 CLKBUF_X1 _34451_ (.A(net182),
    .Z(_16908_));
 CLKBUF_X1 _34452_ (.A(_00833_),
    .Z(_00234_));
 CLKBUF_X1 _34453_ (.A(net181),
    .Z(_16909_));
 CLKBUF_X1 _34454_ (.A(_00834_),
    .Z(_00235_));
 CLKBUF_X1 _34455_ (.A(net180),
    .Z(_16910_));
 CLKBUF_X1 _34456_ (.A(_00835_),
    .Z(_00236_));
 CLKBUF_X1 _34457_ (.A(net179),
    .Z(_16911_));
 CLKBUF_X1 _34458_ (.A(_00836_),
    .Z(_00237_));
 CLKBUF_X1 _34459_ (.A(net178),
    .Z(_16913_));
 CLKBUF_X1 _34460_ (.A(_00838_),
    .Z(_00239_));
 CLKBUF_X1 _34461_ (.A(net177),
    .Z(_16914_));
 CLKBUF_X1 _34462_ (.A(_00839_),
    .Z(_00240_));
 CLKBUF_X1 _34463_ (.A(net176),
    .Z(_16915_));
 CLKBUF_X1 _34464_ (.A(_00840_),
    .Z(_00241_));
 CLKBUF_X1 _34465_ (.A(net175),
    .Z(_16916_));
 CLKBUF_X1 _34466_ (.A(_00841_),
    .Z(_00242_));
 CLKBUF_X1 _34467_ (.A(net174),
    .Z(_16917_));
 CLKBUF_X1 _34468_ (.A(_00842_),
    .Z(_00243_));
 CLKBUF_X1 _34469_ (.A(net173),
    .Z(_16918_));
 CLKBUF_X1 _34470_ (.A(_00843_),
    .Z(_00244_));
 CLKBUF_X1 _34471_ (.A(net172),
    .Z(_16919_));
 CLKBUF_X1 _34472_ (.A(_00844_),
    .Z(_00245_));
 CLKBUF_X1 _34473_ (.A(net171),
    .Z(_16920_));
 CLKBUF_X1 _34474_ (.A(_00845_),
    .Z(_00246_));
 CLKBUF_X1 _34475_ (.A(net170),
    .Z(_16921_));
 CLKBUF_X1 _34476_ (.A(_00846_),
    .Z(_00247_));
 CLKBUF_X1 _34477_ (.A(net169),
    .Z(_16922_));
 CLKBUF_X1 _34478_ (.A(_00847_),
    .Z(_00248_));
 CLKBUF_X1 _34479_ (.A(net168),
    .Z(_16924_));
 CLKBUF_X1 _34480_ (.A(_00849_),
    .Z(_00250_));
 CLKBUF_X1 _34481_ (.A(net167),
    .Z(_16925_));
 CLKBUF_X1 _34482_ (.A(_00850_),
    .Z(_00251_));
 CLKBUF_X1 _34483_ (.A(net166),
    .Z(_16926_));
 CLKBUF_X1 _34484_ (.A(_00851_),
    .Z(_00252_));
 CLKBUF_X1 _34485_ (.A(net165),
    .Z(_16927_));
 CLKBUF_X1 _34486_ (.A(_00852_),
    .Z(_00253_));
 CLKBUF_X1 _34487_ (.A(net164),
    .Z(_16928_));
 CLKBUF_X1 _34488_ (.A(_00853_),
    .Z(_00254_));
 CLKBUF_X1 _34489_ (.A(net163),
    .Z(_16929_));
 CLKBUF_X1 _34490_ (.A(_00854_),
    .Z(_00255_));
 CLKBUF_X1 _34491_ (.A(\sa00[5] ),
    .Z(_16684_));
 CLKBUF_X1 _34492_ (.A(\sa00[4] ),
    .Z(_16683_));
 CLKBUF_X1 _34493_ (.A(\sa00[7] ),
    .Z(_16686_));
 CLKBUF_X1 _34494_ (.A(\sa00[6] ),
    .Z(_16685_));
 CLKBUF_X1 _34495_ (.A(\sa00[1] ),
    .Z(_16680_));
 CLKBUF_X2 _34496_ (.A(\sa00[0] ),
    .Z(_16679_));
 CLKBUF_X2 _34497_ (.A(\sa00[2] ),
    .Z(_16681_));
 CLKBUF_X2 _34498_ (.A(\sa00[3] ),
    .Z(_16682_));
 CLKBUF_X1 _34499_ (.A(\sa11[5] ),
    .Z(_16724_));
 CLKBUF_X1 _34500_ (.A(\sa11[4] ),
    .Z(_16723_));
 CLKBUF_X1 _34501_ (.A(\sa11[7] ),
    .Z(_16726_));
 CLKBUF_X1 _34502_ (.A(\sa11[6] ),
    .Z(_16725_));
 CLKBUF_X2 _34503_ (.A(\sa11[1] ),
    .Z(_16720_));
 BUF_X2 _34504_ (.A(\sa11[0] ),
    .Z(_16719_));
 BUF_X2 _34505_ (.A(\sa11[2] ),
    .Z(_16721_));
 CLKBUF_X2 _34506_ (.A(\sa11[3] ),
    .Z(_16722_));
 CLKBUF_X1 _34507_ (.A(\sa22[5] ),
    .Z(_16764_));
 BUF_X1 _34508_ (.A(\sa22[4] ),
    .Z(_16763_));
 CLKBUF_X1 _34509_ (.A(\sa22[7] ),
    .Z(_16766_));
 CLKBUF_X1 _34510_ (.A(\sa22[6] ),
    .Z(_16765_));
 BUF_X2 _34511_ (.A(\sa22[1] ),
    .Z(_16760_));
 CLKBUF_X2 _34512_ (.A(\sa22[0] ),
    .Z(_16759_));
 BUF_X2 _34513_ (.A(\sa22[2] ),
    .Z(_16761_));
 BUF_X1 _34514_ (.A(\sa22[3] ),
    .Z(_16762_));
 CLKBUF_X2 _34515_ (.A(\sa33[0] ),
    .Z(_16799_));
 CLKBUF_X2 _34516_ (.A(\sa33[1] ),
    .Z(_16800_));
 CLKBUF_X2 _34517_ (.A(\sa33[3] ),
    .Z(_16802_));
 BUF_X2 _34518_ (.A(\sa33[2] ),
    .Z(_16801_));
 CLKBUF_X1 _34519_ (.A(\sa33[5] ),
    .Z(_16804_));
 BUF_X1 _34520_ (.A(\sa33[4] ),
    .Z(_16803_));
 CLKBUF_X1 _34521_ (.A(\sa33[6] ),
    .Z(_16805_));
 CLKBUF_X1 _34522_ (.A(\sa33[7] ),
    .Z(_16806_));
 CLKBUF_X1 _34523_ (.A(\text_in_r[96] ),
    .Z(_17058_));
 CLKBUF_X1 _34524_ (.A(_00700_),
    .Z(_00101_));
 CLKBUF_X1 _34525_ (.A(net162),
    .Z(_16930_));
 CLKBUF_X1 _34526_ (.A(_00855_),
    .Z(_00256_));
 CLKBUF_X1 _34527_ (.A(\text_in_r[97] ),
    .Z(_17059_));
 CLKBUF_X1 _34528_ (.A(net161),
    .Z(_16931_));
 CLKBUF_X1 _34529_ (.A(_00856_),
    .Z(_00257_));
 CLKBUF_X1 _34530_ (.A(\text_in_r[98] ),
    .Z(_17060_));
 CLKBUF_X1 _34531_ (.A(net160),
    .Z(_16932_));
 CLKBUF_X1 _34532_ (.A(_00857_),
    .Z(_00258_));
 CLKBUF_X1 _34533_ (.A(\text_in_r[99] ),
    .Z(_17061_));
 CLKBUF_X1 _34534_ (.A(net159),
    .Z(_16933_));
 CLKBUF_X1 _34535_ (.A(_00858_),
    .Z(_00259_));
 CLKBUF_X1 _34536_ (.A(\text_in_r[100] ),
    .Z(_16936_));
 CLKBUF_X1 _34537_ (.A(net158),
    .Z(_16808_));
 CLKBUF_X1 _34538_ (.A(_00733_),
    .Z(_00134_));
 CLKBUF_X1 _34539_ (.A(\text_in_r[101] ),
    .Z(_16937_));
 CLKBUF_X1 _34540_ (.A(net157),
    .Z(_16809_));
 CLKBUF_X1 _34541_ (.A(_00734_),
    .Z(_00135_));
 CLKBUF_X1 _34542_ (.A(\text_in_r[102] ),
    .Z(_16938_));
 CLKBUF_X1 _34543_ (.A(net156),
    .Z(_16810_));
 CLKBUF_X1 _34544_ (.A(_00735_),
    .Z(_00136_));
 CLKBUF_X1 _34545_ (.A(\text_in_r[103] ),
    .Z(_16939_));
 CLKBUF_X1 _34546_ (.A(net155),
    .Z(_16811_));
 CLKBUF_X1 _34547_ (.A(_00736_),
    .Z(_00137_));
 CLKBUF_X1 _34548_ (.A(\text_in_r[104] ),
    .Z(_16940_));
 CLKBUF_X1 _34549_ (.A(net154),
    .Z(_16812_));
 CLKBUF_X1 _34550_ (.A(_00737_),
    .Z(_00138_));
 CLKBUF_X1 _34551_ (.A(\text_in_r[105] ),
    .Z(_16941_));
 CLKBUF_X1 _34552_ (.A(net153),
    .Z(_16813_));
 CLKBUF_X1 _34553_ (.A(_00738_),
    .Z(_00139_));
 CLKBUF_X1 _34554_ (.A(_00701_),
    .Z(_00102_));
 CLKBUF_X1 _34555_ (.A(\text_in_r[106] ),
    .Z(_16942_));
 CLKBUF_X1 _34556_ (.A(net152),
    .Z(_16814_));
 CLKBUF_X1 _34557_ (.A(_00739_),
    .Z(_00140_));
 CLKBUF_X1 _34558_ (.A(\text_in_r[107] ),
    .Z(_16943_));
 CLKBUF_X1 _34559_ (.A(net151),
    .Z(_16815_));
 CLKBUF_X1 _34560_ (.A(_00740_),
    .Z(_00141_));
 CLKBUF_X1 _34561_ (.A(\text_in_r[108] ),
    .Z(_16944_));
 CLKBUF_X1 _34562_ (.A(net150),
    .Z(_16816_));
 CLKBUF_X1 _34563_ (.A(_00741_),
    .Z(_00142_));
 CLKBUF_X1 _34564_ (.A(\text_in_r[109] ),
    .Z(_16945_));
 CLKBUF_X1 _34565_ (.A(net149),
    .Z(_16817_));
 CLKBUF_X1 _34566_ (.A(_00742_),
    .Z(_00143_));
 CLKBUF_X1 _34567_ (.A(\text_in_r[110] ),
    .Z(_16947_));
 CLKBUF_X1 _34568_ (.A(net148),
    .Z(_16819_));
 CLKBUF_X1 _34569_ (.A(_00744_),
    .Z(_00145_));
 CLKBUF_X1 _34570_ (.A(\text_in_r[111] ),
    .Z(_16948_));
 CLKBUF_X1 _34571_ (.A(net147),
    .Z(_16820_));
 CLKBUF_X1 _34572_ (.A(_00745_),
    .Z(_00146_));
 CLKBUF_X1 _34573_ (.A(\text_in_r[112] ),
    .Z(_16949_));
 CLKBUF_X1 _34574_ (.A(net146),
    .Z(_16821_));
 CLKBUF_X1 _34575_ (.A(_00746_),
    .Z(_00147_));
 CLKBUF_X1 _34576_ (.A(\text_in_r[113] ),
    .Z(_16950_));
 CLKBUF_X1 _34577_ (.A(net145),
    .Z(_16822_));
 CLKBUF_X1 _34578_ (.A(_00747_),
    .Z(_00148_));
 CLKBUF_X1 _34579_ (.A(\text_in_r[114] ),
    .Z(_16951_));
 CLKBUF_X1 _34580_ (.A(net144),
    .Z(_16823_));
 CLKBUF_X1 _34581_ (.A(_00748_),
    .Z(_00149_));
 CLKBUF_X1 _34582_ (.A(\text_in_r[115] ),
    .Z(_16952_));
 CLKBUF_X1 _34583_ (.A(net143),
    .Z(_16824_));
 CLKBUF_X1 _34584_ (.A(_00749_),
    .Z(_00150_));
 CLKBUF_X1 _34585_ (.A(_00702_),
    .Z(_00103_));
 CLKBUF_X1 _34586_ (.A(\text_in_r[116] ),
    .Z(_16953_));
 CLKBUF_X1 _34587_ (.A(net142),
    .Z(_16825_));
 CLKBUF_X1 _34588_ (.A(_00750_),
    .Z(_00151_));
 CLKBUF_X1 _34589_ (.A(\text_in_r[117] ),
    .Z(_16954_));
 CLKBUF_X1 _34590_ (.A(net141),
    .Z(_16826_));
 CLKBUF_X1 _34591_ (.A(_00751_),
    .Z(_00152_));
 CLKBUF_X1 _34592_ (.A(\text_in_r[118] ),
    .Z(_16955_));
 CLKBUF_X1 _34593_ (.A(net140),
    .Z(_16827_));
 CLKBUF_X1 _34594_ (.A(_00752_),
    .Z(_00153_));
 CLKBUF_X1 _34595_ (.A(\text_in_r[119] ),
    .Z(_16956_));
 CLKBUF_X1 _34596_ (.A(net139),
    .Z(_16828_));
 CLKBUF_X1 _34597_ (.A(_00753_),
    .Z(_00154_));
 CLKBUF_X1 _34598_ (.A(\text_in_r[120] ),
    .Z(_16958_));
 CLKBUF_X1 _34599_ (.A(net138),
    .Z(_16830_));
 CLKBUF_X1 _34600_ (.A(_00755_),
    .Z(_00156_));
 CLKBUF_X1 _34601_ (.A(\text_in_r[121] ),
    .Z(_16959_));
 CLKBUF_X1 _34602_ (.A(net137),
    .Z(_16831_));
 CLKBUF_X1 _34603_ (.A(_00756_),
    .Z(_00157_));
 CLKBUF_X1 _34604_ (.A(\text_in_r[122] ),
    .Z(_16960_));
 CLKBUF_X1 _34605_ (.A(net136),
    .Z(_16832_));
 CLKBUF_X1 _34606_ (.A(_00757_),
    .Z(_00158_));
 CLKBUF_X1 _34607_ (.A(\text_in_r[123] ),
    .Z(_16961_));
 CLKBUF_X1 _34608_ (.A(net135),
    .Z(_16833_));
 CLKBUF_X1 _34609_ (.A(_00758_),
    .Z(_00159_));
 CLKBUF_X1 _34610_ (.A(\text_in_r[124] ),
    .Z(_16962_));
 CLKBUF_X1 _34611_ (.A(net134),
    .Z(_16834_));
 CLKBUF_X1 _34612_ (.A(_00759_),
    .Z(_00160_));
 CLKBUF_X1 _34613_ (.A(\text_in_r[125] ),
    .Z(_16963_));
 CLKBUF_X1 _34614_ (.A(net133),
    .Z(_16835_));
 CLKBUF_X1 _34615_ (.A(_00760_),
    .Z(_00161_));
 CLKBUF_X1 _34616_ (.A(_00703_),
    .Z(_00104_));
 CLKBUF_X1 _34617_ (.A(\text_in_r[126] ),
    .Z(_16964_));
 CLKBUF_X1 _34618_ (.A(net132),
    .Z(_16836_));
 CLKBUF_X1 _34619_ (.A(_00761_),
    .Z(_00162_));
 CLKBUF_X1 _34620_ (.A(\text_in_r[127] ),
    .Z(_16965_));
 CLKBUF_X1 _34621_ (.A(net131),
    .Z(_16837_));
 CLKBUF_X1 _34622_ (.A(_00762_),
    .Z(_00163_));
 CLKBUF_X1 _34623_ (.A(_00704_),
    .Z(_00105_));
 CLKBUF_X1 _34624_ (.A(_00705_),
    .Z(_00106_));
 CLKBUF_X1 _34625_ (.A(_00706_),
    .Z(_00107_));
 CLKBUF_X1 _34626_ (.A(_00707_),
    .Z(_00108_));
 CLKBUF_X1 _34627_ (.A(_00668_),
    .Z(_00069_));
 CLKBUF_X1 _34628_ (.A(_00669_),
    .Z(_00070_));
 CLKBUF_X1 _34629_ (.A(_00670_),
    .Z(_00071_));
 CLKBUF_X1 _34630_ (.A(_00671_),
    .Z(_00072_));
 CLKBUF_X1 _34631_ (.A(_00672_),
    .Z(_00073_));
 CLKBUF_X1 _34632_ (.A(_00673_),
    .Z(_00074_));
 CLKBUF_X1 _34633_ (.A(_00674_),
    .Z(_00075_));
 CLKBUF_X1 _34634_ (.A(_00675_),
    .Z(_00076_));
 CLKBUF_X1 _34635_ (.A(_00636_),
    .Z(_00037_));
 CLKBUF_X1 _34636_ (.A(_00637_),
    .Z(_00038_));
 CLKBUF_X1 _34637_ (.A(_00638_),
    .Z(_00039_));
 CLKBUF_X1 _34638_ (.A(_00639_),
    .Z(_00040_));
 CLKBUF_X1 _34639_ (.A(_00640_),
    .Z(_00041_));
 CLKBUF_X1 _34640_ (.A(_00641_),
    .Z(_00042_));
 CLKBUF_X1 _34641_ (.A(_00642_),
    .Z(_00043_));
 CLKBUF_X1 _34642_ (.A(_00643_),
    .Z(_00044_));
 CLKBUF_X1 _34643_ (.A(_00604_),
    .Z(_00005_));
 CLKBUF_X1 _34644_ (.A(_00605_),
    .Z(_00006_));
 CLKBUF_X1 _34645_ (.A(_00606_),
    .Z(_00007_));
 CLKBUF_X1 _34646_ (.A(_00607_),
    .Z(_00008_));
 CLKBUF_X1 _34647_ (.A(_00608_),
    .Z(_00009_));
 CLKBUF_X1 _34648_ (.A(_00609_),
    .Z(_00010_));
 CLKBUF_X1 _34649_ (.A(_00610_),
    .Z(_00011_));
 CLKBUF_X1 _34650_ (.A(_00611_),
    .Z(_00012_));
 CLKBUF_X1 _34651_ (.A(_00603_),
    .Z(_00004_));
 CLKBUF_X1 _34652_ (.A(_00884_),
    .Z(_00285_));
 CLKBUF_X1 _34653_ (.A(_00885_),
    .Z(_00286_));
 CLKBUF_X1 _34654_ (.A(_00886_),
    .Z(_00287_));
 CLKBUF_X1 _34655_ (.A(_00887_),
    .Z(_00288_));
 CLKBUF_X1 _34656_ (.A(_00888_),
    .Z(_00289_));
 CLKBUF_X1 _34657_ (.A(_00889_),
    .Z(_00290_));
 CLKBUF_X1 _34658_ (.A(_00890_),
    .Z(_00291_));
 CLKBUF_X1 _34659_ (.A(_00891_),
    .Z(_00292_));
 CLKBUF_X1 _34660_ (.A(_00980_),
    .Z(_00381_));
 CLKBUF_X1 _34661_ (.A(_00981_),
    .Z(_00382_));
 CLKBUF_X1 _34662_ (.A(_00982_),
    .Z(_00383_));
 CLKBUF_X1 _34663_ (.A(_00983_),
    .Z(_00384_));
 CLKBUF_X1 _34664_ (.A(_00984_),
    .Z(_00385_));
 CLKBUF_X1 _34665_ (.A(_00985_),
    .Z(_00386_));
 CLKBUF_X1 _34666_ (.A(_00986_),
    .Z(_00387_));
 CLKBUF_X1 _34667_ (.A(_00987_),
    .Z(_00388_));
 CLKBUF_X1 _34668_ (.A(_00940_),
    .Z(_00341_));
 CLKBUF_X1 _34669_ (.A(_00941_),
    .Z(_00342_));
 CLKBUF_X1 _34670_ (.A(_00942_),
    .Z(_00343_));
 CLKBUF_X1 _34671_ (.A(_00943_),
    .Z(_00344_));
 CLKBUF_X1 _34672_ (.A(_00944_),
    .Z(_00345_));
 CLKBUF_X1 _34673_ (.A(_00945_),
    .Z(_00346_));
 CLKBUF_X1 _34674_ (.A(_00946_),
    .Z(_00347_));
 CLKBUF_X1 _34675_ (.A(_00947_),
    .Z(_00348_));
 CLKBUF_X1 _34676_ (.A(_00908_),
    .Z(_00309_));
 CLKBUF_X1 _34677_ (.A(_00909_),
    .Z(_00310_));
 CLKBUF_X1 _34678_ (.A(_00910_),
    .Z(_00311_));
 CLKBUF_X1 _34679_ (.A(_00911_),
    .Z(_00312_));
 CLKBUF_X1 _34680_ (.A(_00912_),
    .Z(_00313_));
 CLKBUF_X1 _34681_ (.A(_00913_),
    .Z(_00314_));
 CLKBUF_X1 _34682_ (.A(_00914_),
    .Z(_00315_));
 CLKBUF_X1 _34683_ (.A(_00915_),
    .Z(_00316_));
 CLKBUF_X1 _34684_ (.A(_00876_),
    .Z(_00277_));
 CLKBUF_X1 _34685_ (.A(_00877_),
    .Z(_00278_));
 CLKBUF_X1 _34686_ (.A(_00878_),
    .Z(_00279_));
 CLKBUF_X1 _34687_ (.A(_00879_),
    .Z(_00280_));
 CLKBUF_X1 _34688_ (.A(_00880_),
    .Z(_00281_));
 CLKBUF_X1 _34689_ (.A(_00881_),
    .Z(_00282_));
 CLKBUF_X1 _34690_ (.A(_00882_),
    .Z(_00283_));
 CLKBUF_X1 _34691_ (.A(_00883_),
    .Z(_00284_));
 CLKBUF_X1 _34692_ (.A(_00972_),
    .Z(_00373_));
 CLKBUF_X1 _34693_ (.A(_00973_),
    .Z(_00374_));
 CLKBUF_X1 _34694_ (.A(_00974_),
    .Z(_00375_));
 CLKBUF_X1 _34695_ (.A(_00975_),
    .Z(_00376_));
 CLKBUF_X1 _34696_ (.A(_00976_),
    .Z(_00377_));
 CLKBUF_X1 _34697_ (.A(_00977_),
    .Z(_00378_));
 CLKBUF_X1 _34698_ (.A(_00978_),
    .Z(_00379_));
 CLKBUF_X1 _34699_ (.A(_00979_),
    .Z(_00380_));
 CLKBUF_X1 _34700_ (.A(_00932_),
    .Z(_00333_));
 CLKBUF_X1 _34701_ (.A(_00933_),
    .Z(_00334_));
 CLKBUF_X1 _34702_ (.A(_00934_),
    .Z(_00335_));
 CLKBUF_X1 _34703_ (.A(_00935_),
    .Z(_00336_));
 CLKBUF_X1 _34704_ (.A(_00936_),
    .Z(_00337_));
 CLKBUF_X1 _34705_ (.A(_00937_),
    .Z(_00338_));
 CLKBUF_X1 _34706_ (.A(_00938_),
    .Z(_00339_));
 CLKBUF_X1 _34707_ (.A(_00939_),
    .Z(_00340_));
 CLKBUF_X1 _34708_ (.A(_00900_),
    .Z(_00301_));
 CLKBUF_X1 _34709_ (.A(_00901_),
    .Z(_00302_));
 CLKBUF_X1 _34710_ (.A(_00902_),
    .Z(_00303_));
 CLKBUF_X1 _34711_ (.A(_00903_),
    .Z(_00304_));
 CLKBUF_X1 _34712_ (.A(_00904_),
    .Z(_00305_));
 CLKBUF_X1 _34713_ (.A(_00905_),
    .Z(_00306_));
 CLKBUF_X1 _34714_ (.A(_00906_),
    .Z(_00307_));
 CLKBUF_X1 _34715_ (.A(_00907_),
    .Z(_00308_));
 CLKBUF_X1 _34716_ (.A(_00868_),
    .Z(_00269_));
 CLKBUF_X1 _34717_ (.A(_00869_),
    .Z(_00270_));
 CLKBUF_X1 _34718_ (.A(_00870_),
    .Z(_00271_));
 CLKBUF_X1 _34719_ (.A(_00871_),
    .Z(_00272_));
 CLKBUF_X1 _34720_ (.A(_00872_),
    .Z(_00273_));
 CLKBUF_X1 _34721_ (.A(_00873_),
    .Z(_00274_));
 CLKBUF_X1 _34722_ (.A(_00874_),
    .Z(_00275_));
 CLKBUF_X1 _34723_ (.A(_00875_),
    .Z(_00276_));
 CLKBUF_X1 _34724_ (.A(_00956_),
    .Z(_00357_));
 CLKBUF_X1 _34725_ (.A(_00957_),
    .Z(_00358_));
 CLKBUF_X1 _34726_ (.A(_00958_),
    .Z(_00359_));
 CLKBUF_X1 _34727_ (.A(_00959_),
    .Z(_00360_));
 CLKBUF_X1 _34728_ (.A(_00960_),
    .Z(_00361_));
 CLKBUF_X1 _34729_ (.A(_00961_),
    .Z(_00362_));
 CLKBUF_X1 _34730_ (.A(_00962_),
    .Z(_00363_));
 CLKBUF_X1 _34731_ (.A(_00963_),
    .Z(_00364_));
 CLKBUF_X1 _34732_ (.A(_00924_),
    .Z(_00325_));
 CLKBUF_X1 _34733_ (.A(_00925_),
    .Z(_00326_));
 CLKBUF_X1 _34734_ (.A(_00926_),
    .Z(_00327_));
 CLKBUF_X1 _34735_ (.A(_00927_),
    .Z(_00328_));
 CLKBUF_X1 _34736_ (.A(_00928_),
    .Z(_00329_));
 CLKBUF_X1 _34737_ (.A(_00929_),
    .Z(_00330_));
 CLKBUF_X1 _34738_ (.A(_00930_),
    .Z(_00331_));
 CLKBUF_X1 _34739_ (.A(_00931_),
    .Z(_00332_));
 CLKBUF_X1 _34740_ (.A(_00892_),
    .Z(_00293_));
 CLKBUF_X1 _34741_ (.A(_00893_),
    .Z(_00294_));
 CLKBUF_X1 _34742_ (.A(_00894_),
    .Z(_00295_));
 CLKBUF_X1 _34743_ (.A(_00895_),
    .Z(_00296_));
 CLKBUF_X1 _34744_ (.A(_00896_),
    .Z(_00297_));
 CLKBUF_X1 _34745_ (.A(_00897_),
    .Z(_00298_));
 CLKBUF_X1 _34746_ (.A(_00898_),
    .Z(_00299_));
 CLKBUF_X1 _34747_ (.A(_00899_),
    .Z(_00300_));
 CLKBUF_X1 _34748_ (.A(_00860_),
    .Z(_00261_));
 CLKBUF_X1 _34749_ (.A(_00861_),
    .Z(_00262_));
 CLKBUF_X1 _34750_ (.A(_00862_),
    .Z(_00263_));
 CLKBUF_X1 _34751_ (.A(_00863_),
    .Z(_00264_));
 CLKBUF_X1 _34752_ (.A(_00864_),
    .Z(_00265_));
 CLKBUF_X1 _34753_ (.A(_00865_),
    .Z(_00266_));
 CLKBUF_X1 _34754_ (.A(_00866_),
    .Z(_00267_));
 CLKBUF_X1 _34755_ (.A(_00867_),
    .Z(_00268_));
 CLKBUF_X1 _34756_ (.A(_00948_),
    .Z(_00349_));
 CLKBUF_X1 _34757_ (.A(_00949_),
    .Z(_00350_));
 CLKBUF_X1 _34758_ (.A(_00950_),
    .Z(_00351_));
 CLKBUF_X1 _34759_ (.A(_00951_),
    .Z(_00352_));
 CLKBUF_X1 _34760_ (.A(_00952_),
    .Z(_00353_));
 CLKBUF_X1 _34761_ (.A(_00953_),
    .Z(_00354_));
 CLKBUF_X1 _34762_ (.A(_00954_),
    .Z(_00355_));
 CLKBUF_X1 _34763_ (.A(_00955_),
    .Z(_00356_));
 CLKBUF_X1 _34764_ (.A(_00916_),
    .Z(_00317_));
 CLKBUF_X1 _34765_ (.A(_00917_),
    .Z(_00318_));
 CLKBUF_X1 _34766_ (.A(_00918_),
    .Z(_00319_));
 CLKBUF_X1 _34767_ (.A(_00919_),
    .Z(_00320_));
 CLKBUF_X1 _34768_ (.A(_00920_),
    .Z(_00321_));
 CLKBUF_X1 _34769_ (.A(_00921_),
    .Z(_00322_));
 CLKBUF_X1 _34770_ (.A(_00922_),
    .Z(_00323_));
 CLKBUF_X1 _34771_ (.A(_00923_),
    .Z(_00324_));
 CLKBUF_X1 _34772_ (.A(_00964_),
    .Z(_00365_));
 CLKBUF_X1 _34773_ (.A(_00965_),
    .Z(_00366_));
 CLKBUF_X1 _34774_ (.A(_00966_),
    .Z(_00367_));
 CLKBUF_X1 _34775_ (.A(_00967_),
    .Z(_00368_));
 CLKBUF_X1 _34776_ (.A(_00968_),
    .Z(_00369_));
 CLKBUF_X1 _34777_ (.A(_00969_),
    .Z(_00370_));
 CLKBUF_X1 _34778_ (.A(_00970_),
    .Z(_00371_));
 CLKBUF_X1 _34779_ (.A(_00971_),
    .Z(_00372_));
 DFF_X1 _34780_ (.D(_00595_),
    .CK(clk),
    .Q(\u0.r0.rcnt[0] ),
    .QN(_17195_));
 DFF_X1 _34781_ (.D(_00596_),
    .CK(clk),
    .Q(\u0.r0.rcnt[1] ),
    .QN(_17196_));
 DFF_X1 _34782_ (.D(_00597_),
    .CK(clk),
    .Q(\u0.r0.rcnt[2] ),
    .QN(_17197_));
 DFF_X1 _34783_ (.D(_00598_),
    .CK(clk),
    .Q(\u0.r0.rcnt[3] ),
    .QN(_17198_));
 DFF_X1 _34784_ (.D(_00587_),
    .CK(clk),
    .Q(\u0.r0.out[24] ),
    .QN(_00414_));
 DFF_X1 _34785_ (.D(_00588_),
    .CK(clk),
    .Q(\u0.r0.out[25] ),
    .QN(_00416_));
 DFF_X1 _34786_ (.D(_00589_),
    .CK(clk),
    .Q(\u0.r0.out[26] ),
    .QN(_00418_));
 DFF_X1 _34787_ (.D(_00590_),
    .CK(clk),
    .Q(\u0.r0.out[27] ),
    .QN(_00420_));
 DFF_X1 _34788_ (.D(_00591_),
    .CK(clk),
    .Q(\u0.r0.out[28] ),
    .QN(_00422_));
 DFF_X1 _34789_ (.D(_00592_),
    .CK(clk),
    .Q(\u0.r0.out[29] ),
    .QN(_00424_));
 DFF_X1 _34790_ (.D(_00593_),
    .CK(clk),
    .Q(\u0.r0.out[30] ),
    .QN(_00426_));
 DFF_X1 _34791_ (.D(_00594_),
    .CK(clk),
    .Q(\u0.r0.out[31] ),
    .QN(_00428_));
 DFF_X1 _34792_ (.D(_00555_),
    .CK(clk),
    .Q(\u0.tmp_w[0] ),
    .QN(_17199_));
 DFF_X1 _34793_ (.D(_00566_),
    .CK(clk),
    .Q(\u0.tmp_w[1] ),
    .QN(_17200_));
 DFF_X1 _34794_ (.D(_00577_),
    .CK(clk),
    .Q(\u0.tmp_w[2] ),
    .QN(_17201_));
 DFF_X1 _34795_ (.D(_00580_),
    .CK(clk),
    .Q(\u0.tmp_w[3] ),
    .QN(_17202_));
 DFF_X1 _34796_ (.D(_00581_),
    .CK(clk),
    .Q(\u0.tmp_w[4] ),
    .QN(_17203_));
 DFF_X1 _34797_ (.D(_00582_),
    .CK(clk),
    .Q(\u0.tmp_w[5] ),
    .QN(_17204_));
 DFF_X1 _34798_ (.D(_00583_),
    .CK(clk),
    .Q(\u0.tmp_w[6] ),
    .QN(_17205_));
 DFF_X1 _34799_ (.D(_00584_),
    .CK(clk),
    .Q(\u0.tmp_w[7] ),
    .QN(_17206_));
 DFF_X1 _34800_ (.D(_00585_),
    .CK(clk),
    .Q(\u0.tmp_w[8] ),
    .QN(_00450_));
 DFF_X1 _34801_ (.D(_00586_),
    .CK(clk),
    .Q(\u0.tmp_w[9] ),
    .QN(_17207_));
 DFF_X1 _34802_ (.D(_00556_),
    .CK(clk),
    .Q(\u0.tmp_w[10] ),
    .QN(_17208_));
 DFF_X1 _34803_ (.D(_00557_),
    .CK(clk),
    .Q(\u0.tmp_w[11] ),
    .QN(_17209_));
 DFF_X1 _34804_ (.D(_00558_),
    .CK(clk),
    .Q(\u0.tmp_w[12] ),
    .QN(_17210_));
 DFF_X1 _34805_ (.D(_00559_),
    .CK(clk),
    .Q(\u0.tmp_w[13] ),
    .QN(_17211_));
 DFF_X1 _34806_ (.D(_00560_),
    .CK(clk),
    .Q(\u0.tmp_w[14] ),
    .QN(_17212_));
 DFF_X1 _34807_ (.D(_00561_),
    .CK(clk),
    .Q(\u0.tmp_w[15] ),
    .QN(_17213_));
 DFF_X1 _34808_ (.D(_00562_),
    .CK(clk),
    .Q(\u0.tmp_w[16] ),
    .QN(_00451_));
 DFF_X1 _34809_ (.D(_00563_),
    .CK(clk),
    .Q(\u0.tmp_w[17] ),
    .QN(_00452_));
 DFF_X1 _34810_ (.D(_00564_),
    .CK(clk),
    .Q(\u0.tmp_w[18] ),
    .QN(_17214_));
 DFF_X1 _34811_ (.D(_00565_),
    .CK(clk),
    .Q(\u0.tmp_w[19] ),
    .QN(_17215_));
 DFF_X1 _34812_ (.D(_00567_),
    .CK(clk),
    .Q(\u0.tmp_w[20] ),
    .QN(_17216_));
 DFF_X1 _34813_ (.D(_00568_),
    .CK(clk),
    .Q(\u0.tmp_w[21] ),
    .QN(_00453_));
 DFF_X1 _34814_ (.D(_00569_),
    .CK(clk),
    .Q(\u0.tmp_w[22] ),
    .QN(_00454_));
 DFF_X1 _34815_ (.D(_00570_),
    .CK(clk),
    .Q(\u0.tmp_w[23] ),
    .QN(_17217_));
 DFF_X1 _34816_ (.D(_00571_),
    .CK(clk),
    .Q(\u0.tmp_w[24] ),
    .QN(_00455_));
 DFF_X1 _34817_ (.D(_00572_),
    .CK(clk),
    .Q(\u0.tmp_w[25] ),
    .QN(_00456_));
 DFF_X1 _34818_ (.D(_00573_),
    .CK(clk),
    .Q(\u0.tmp_w[26] ),
    .QN(_17218_));
 DFF_X1 _34819_ (.D(_00574_),
    .CK(clk),
    .Q(\u0.tmp_w[27] ),
    .QN(_17219_));
 DFF_X1 _34820_ (.D(_00575_),
    .CK(clk),
    .Q(\u0.tmp_w[28] ),
    .QN(_17220_));
 DFF_X1 _34821_ (.D(_00576_),
    .CK(clk),
    .Q(\u0.tmp_w[29] ),
    .QN(_00457_));
 DFF_X1 _34822_ (.D(_00578_),
    .CK(clk),
    .Q(\u0.tmp_w[30] ),
    .QN(_00458_));
 DFF_X1 _34823_ (.D(_00579_),
    .CK(clk),
    .Q(\u0.tmp_w[31] ),
    .QN(_17221_));
 DFF_X1 _34824_ (.D(_00000_),
    .CK(clk),
    .Q(\dcnt[0] ),
    .QN(_17222_));
 DFF_X1 _34825_ (.D(_00001_),
    .CK(clk),
    .Q(\dcnt[1] ),
    .QN(_00446_));
 DFF_X1 _34826_ (.D(_00002_),
    .CK(clk),
    .Q(\dcnt[2] ),
    .QN(_00447_));
 DFF_X1 _34827_ (.D(_00003_),
    .CK(clk),
    .Q(\dcnt[3] ),
    .QN(_00448_));
 DFF_X1 _34828_ (.D(_00004_),
    .CK(clk),
    .Q(net259),
    .QN(_17223_));
 DFF_X1 _34829_ (.D(_00133_),
    .CK(clk),
    .Q(\text_in_r[0] ),
    .QN(_17224_));
 DFF_X1 _34830_ (.D(_00172_),
    .CK(clk),
    .Q(\text_in_r[1] ),
    .QN(_17225_));
 DFF_X1 _34831_ (.D(_00183_),
    .CK(clk),
    .Q(\text_in_r[2] ),
    .QN(_17226_));
 DFF_X1 _34832_ (.D(_00194_),
    .CK(clk),
    .Q(\text_in_r[3] ),
    .QN(_17227_));
 DFF_X1 _34833_ (.D(_00205_),
    .CK(clk),
    .Q(\text_in_r[4] ),
    .QN(_17228_));
 DFF_X1 _34834_ (.D(_00216_),
    .CK(clk),
    .Q(\text_in_r[5] ),
    .QN(_17229_));
 DFF_X1 _34835_ (.D(_00227_),
    .CK(clk),
    .Q(\text_in_r[6] ),
    .QN(_17230_));
 DFF_X1 _34836_ (.D(_00238_),
    .CK(clk),
    .Q(\text_in_r[7] ),
    .QN(_17231_));
 DFF_X1 _34837_ (.D(_00249_),
    .CK(clk),
    .Q(\text_in_r[8] ),
    .QN(_17232_));
 DFF_X1 _34838_ (.D(_00260_),
    .CK(clk),
    .Q(\text_in_r[9] ),
    .QN(_17233_));
 DFF_X1 _34839_ (.D(_00144_),
    .CK(clk),
    .Q(\text_in_r[10] ),
    .QN(_17234_));
 DFF_X1 _34840_ (.D(_00155_),
    .CK(clk),
    .Q(\text_in_r[11] ),
    .QN(_17235_));
 DFF_X1 _34841_ (.D(_00164_),
    .CK(clk),
    .Q(\text_in_r[12] ),
    .QN(_17236_));
 DFF_X1 _34842_ (.D(_00165_),
    .CK(clk),
    .Q(\text_in_r[13] ),
    .QN(_17237_));
 DFF_X1 _34843_ (.D(_00166_),
    .CK(clk),
    .Q(\text_in_r[14] ),
    .QN(_17238_));
 DFF_X1 _34844_ (.D(_00167_),
    .CK(clk),
    .Q(\text_in_r[15] ),
    .QN(_17239_));
 DFF_X1 _34845_ (.D(_00168_),
    .CK(clk),
    .Q(\text_in_r[16] ),
    .QN(_17240_));
 DFF_X1 _34846_ (.D(_00169_),
    .CK(clk),
    .Q(\text_in_r[17] ),
    .QN(_17241_));
 DFF_X1 _34847_ (.D(_00170_),
    .CK(clk),
    .Q(\text_in_r[18] ),
    .QN(_17242_));
 DFF_X1 _34848_ (.D(_00171_),
    .CK(clk),
    .Q(\text_in_r[19] ),
    .QN(_17243_));
 DFF_X1 _34849_ (.D(_00173_),
    .CK(clk),
    .Q(\text_in_r[20] ),
    .QN(_17244_));
 DFF_X1 _34850_ (.D(_00174_),
    .CK(clk),
    .Q(\text_in_r[21] ),
    .QN(_17245_));
 DFF_X1 _34851_ (.D(_00175_),
    .CK(clk),
    .Q(\text_in_r[22] ),
    .QN(_17246_));
 DFF_X1 _34852_ (.D(_00176_),
    .CK(clk),
    .Q(\text_in_r[23] ),
    .QN(_17247_));
 DFF_X1 _34853_ (.D(_00177_),
    .CK(clk),
    .Q(\text_in_r[24] ),
    .QN(_17248_));
 DFF_X1 _34854_ (.D(_00178_),
    .CK(clk),
    .Q(\text_in_r[25] ),
    .QN(_17249_));
 DFF_X1 _34855_ (.D(_00179_),
    .CK(clk),
    .Q(\text_in_r[26] ),
    .QN(_17250_));
 DFF_X1 _34856_ (.D(_00180_),
    .CK(clk),
    .Q(\text_in_r[27] ),
    .QN(_17251_));
 DFF_X1 _34857_ (.D(_00181_),
    .CK(clk),
    .Q(\text_in_r[28] ),
    .QN(_17252_));
 DFF_X1 _34858_ (.D(_00182_),
    .CK(clk),
    .Q(\text_in_r[29] ),
    .QN(_17253_));
 DFF_X1 _34859_ (.D(_00184_),
    .CK(clk),
    .Q(\text_in_r[30] ),
    .QN(_17254_));
 DFF_X1 _34860_ (.D(_00185_),
    .CK(clk),
    .Q(\text_in_r[31] ),
    .QN(_17255_));
 DFF_X1 _34861_ (.D(_00186_),
    .CK(clk),
    .Q(\text_in_r[32] ),
    .QN(_17256_));
 DFF_X1 _34862_ (.D(_00187_),
    .CK(clk),
    .Q(\text_in_r[33] ),
    .QN(_17257_));
 DFF_X1 _34863_ (.D(_00188_),
    .CK(clk),
    .Q(\text_in_r[34] ),
    .QN(_17258_));
 DFF_X1 _34864_ (.D(_00189_),
    .CK(clk),
    .Q(\text_in_r[35] ),
    .QN(_17259_));
 DFF_X1 _34865_ (.D(_00190_),
    .CK(clk),
    .Q(\text_in_r[36] ),
    .QN(_17260_));
 DFF_X1 _34866_ (.D(_00191_),
    .CK(clk),
    .Q(\text_in_r[37] ),
    .QN(_17261_));
 DFF_X1 _34867_ (.D(_00192_),
    .CK(clk),
    .Q(\text_in_r[38] ),
    .QN(_17262_));
 DFF_X1 _34868_ (.D(_00193_),
    .CK(clk),
    .Q(\text_in_r[39] ),
    .QN(_17263_));
 DFF_X1 _34869_ (.D(_00195_),
    .CK(clk),
    .Q(\text_in_r[40] ),
    .QN(_17264_));
 DFF_X1 _34870_ (.D(_00196_),
    .CK(clk),
    .Q(\text_in_r[41] ),
    .QN(_17265_));
 DFF_X1 _34871_ (.D(_00197_),
    .CK(clk),
    .Q(\text_in_r[42] ),
    .QN(_17266_));
 DFF_X1 _34872_ (.D(_00198_),
    .CK(clk),
    .Q(\text_in_r[43] ),
    .QN(_17267_));
 DFF_X1 _34873_ (.D(_00199_),
    .CK(clk),
    .Q(\text_in_r[44] ),
    .QN(_17268_));
 DFF_X1 _34874_ (.D(_00200_),
    .CK(clk),
    .Q(\text_in_r[45] ),
    .QN(_17269_));
 DFF_X1 _34875_ (.D(_00201_),
    .CK(clk),
    .Q(\text_in_r[46] ),
    .QN(_17270_));
 DFF_X1 _34876_ (.D(_00202_),
    .CK(clk),
    .Q(\text_in_r[47] ),
    .QN(_17271_));
 DFF_X1 _34877_ (.D(_00203_),
    .CK(clk),
    .Q(\text_in_r[48] ),
    .QN(_17272_));
 DFF_X1 _34878_ (.D(_00204_),
    .CK(clk),
    .Q(\text_in_r[49] ),
    .QN(_17273_));
 DFF_X1 _34879_ (.D(_00206_),
    .CK(clk),
    .Q(\text_in_r[50] ),
    .QN(_17274_));
 DFF_X1 _34880_ (.D(_00207_),
    .CK(clk),
    .Q(\text_in_r[51] ),
    .QN(_17275_));
 DFF_X1 _34881_ (.D(_00208_),
    .CK(clk),
    .Q(\text_in_r[52] ),
    .QN(_17276_));
 DFF_X1 _34882_ (.D(_00209_),
    .CK(clk),
    .Q(\text_in_r[53] ),
    .QN(_17277_));
 DFF_X1 _34883_ (.D(_00210_),
    .CK(clk),
    .Q(\text_in_r[54] ),
    .QN(_17278_));
 DFF_X1 _34884_ (.D(_00211_),
    .CK(clk),
    .Q(\text_in_r[55] ),
    .QN(_17279_));
 DFF_X1 _34885_ (.D(_00212_),
    .CK(clk),
    .Q(\text_in_r[56] ),
    .QN(_17280_));
 DFF_X1 _34886_ (.D(_00213_),
    .CK(clk),
    .Q(\text_in_r[57] ),
    .QN(_17281_));
 DFF_X1 _34887_ (.D(_00214_),
    .CK(clk),
    .Q(\text_in_r[58] ),
    .QN(_17282_));
 DFF_X1 _34888_ (.D(_00215_),
    .CK(clk),
    .Q(\text_in_r[59] ),
    .QN(_17283_));
 DFF_X1 _34889_ (.D(_00217_),
    .CK(clk),
    .Q(\text_in_r[60] ),
    .QN(_17284_));
 DFF_X1 _34890_ (.D(_00218_),
    .CK(clk),
    .Q(\text_in_r[61] ),
    .QN(_17285_));
 DFF_X1 _34891_ (.D(_00219_),
    .CK(clk),
    .Q(\text_in_r[62] ),
    .QN(_17286_));
 DFF_X1 _34892_ (.D(_00220_),
    .CK(clk),
    .Q(\text_in_r[63] ),
    .QN(_17287_));
 DFF_X1 _34893_ (.D(_00221_),
    .CK(clk),
    .Q(\text_in_r[64] ),
    .QN(_17288_));
 DFF_X1 _34894_ (.D(_00222_),
    .CK(clk),
    .Q(\text_in_r[65] ),
    .QN(_17289_));
 DFF_X1 _34895_ (.D(_00223_),
    .CK(clk),
    .Q(\text_in_r[66] ),
    .QN(_17290_));
 DFF_X1 _34896_ (.D(_00224_),
    .CK(clk),
    .Q(\text_in_r[67] ),
    .QN(_17291_));
 DFF_X1 _34897_ (.D(_00225_),
    .CK(clk),
    .Q(\text_in_r[68] ),
    .QN(_17292_));
 DFF_X1 _34898_ (.D(_00226_),
    .CK(clk),
    .Q(\text_in_r[69] ),
    .QN(_17293_));
 DFF_X1 _34899_ (.D(_00228_),
    .CK(clk),
    .Q(\text_in_r[70] ),
    .QN(_17294_));
 DFF_X1 _34900_ (.D(_00229_),
    .CK(clk),
    .Q(\text_in_r[71] ),
    .QN(_17295_));
 DFF_X1 _34901_ (.D(_00230_),
    .CK(clk),
    .Q(\text_in_r[72] ),
    .QN(_17296_));
 DFF_X1 _34902_ (.D(_00231_),
    .CK(clk),
    .Q(\text_in_r[73] ),
    .QN(_17297_));
 DFF_X1 _34903_ (.D(_00232_),
    .CK(clk),
    .Q(\text_in_r[74] ),
    .QN(_17298_));
 DFF_X1 _34904_ (.D(_00233_),
    .CK(clk),
    .Q(\text_in_r[75] ),
    .QN(_17299_));
 DFF_X1 _34905_ (.D(_00234_),
    .CK(clk),
    .Q(\text_in_r[76] ),
    .QN(_17300_));
 DFF_X1 _34906_ (.D(_00235_),
    .CK(clk),
    .Q(\text_in_r[77] ),
    .QN(_17301_));
 DFF_X1 _34907_ (.D(_00236_),
    .CK(clk),
    .Q(\text_in_r[78] ),
    .QN(_17302_));
 DFF_X1 _34908_ (.D(_00237_),
    .CK(clk),
    .Q(\text_in_r[79] ),
    .QN(_17303_));
 DFF_X1 _34909_ (.D(_00239_),
    .CK(clk),
    .Q(\text_in_r[80] ),
    .QN(_17304_));
 DFF_X1 _34910_ (.D(_00240_),
    .CK(clk),
    .Q(\text_in_r[81] ),
    .QN(_17305_));
 DFF_X1 _34911_ (.D(_00241_),
    .CK(clk),
    .Q(\text_in_r[82] ),
    .QN(_17306_));
 DFF_X1 _34912_ (.D(_00242_),
    .CK(clk),
    .Q(\text_in_r[83] ),
    .QN(_17307_));
 DFF_X1 _34913_ (.D(_00243_),
    .CK(clk),
    .Q(\text_in_r[84] ),
    .QN(_17308_));
 DFF_X1 _34914_ (.D(_00244_),
    .CK(clk),
    .Q(\text_in_r[85] ),
    .QN(_17309_));
 DFF_X1 _34915_ (.D(_00245_),
    .CK(clk),
    .Q(\text_in_r[86] ),
    .QN(_17310_));
 DFF_X1 _34916_ (.D(_00246_),
    .CK(clk),
    .Q(\text_in_r[87] ),
    .QN(_17311_));
 DFF_X1 _34917_ (.D(_00247_),
    .CK(clk),
    .Q(\text_in_r[88] ),
    .QN(_17312_));
 DFF_X1 _34918_ (.D(_00248_),
    .CK(clk),
    .Q(\text_in_r[89] ),
    .QN(_17313_));
 DFF_X1 _34919_ (.D(_00250_),
    .CK(clk),
    .Q(\text_in_r[90] ),
    .QN(_17314_));
 DFF_X1 _34920_ (.D(_00251_),
    .CK(clk),
    .Q(\text_in_r[91] ),
    .QN(_17315_));
 DFF_X1 _34921_ (.D(_00252_),
    .CK(clk),
    .Q(\text_in_r[92] ),
    .QN(_17316_));
 DFF_X1 _34922_ (.D(_00253_),
    .CK(clk),
    .Q(\text_in_r[93] ),
    .QN(_17317_));
 DFF_X1 _34923_ (.D(_00254_),
    .CK(clk),
    .Q(\text_in_r[94] ),
    .QN(_17318_));
 DFF_X1 _34924_ (.D(_00255_),
    .CK(clk),
    .Q(\text_in_r[95] ),
    .QN(_17319_));
 DFF_X1 _34925_ (.D(_00256_),
    .CK(clk),
    .Q(\text_in_r[96] ),
    .QN(_17320_));
 DFF_X1 _34926_ (.D(_00257_),
    .CK(clk),
    .Q(\text_in_r[97] ),
    .QN(_17321_));
 DFF_X1 _34927_ (.D(_00258_),
    .CK(clk),
    .Q(\text_in_r[98] ),
    .QN(_17322_));
 DFF_X1 _34928_ (.D(_00259_),
    .CK(clk),
    .Q(\text_in_r[99] ),
    .QN(_17323_));
 DFF_X1 _34929_ (.D(_00134_),
    .CK(clk),
    .Q(\text_in_r[100] ),
    .QN(_17324_));
 DFF_X1 _34930_ (.D(_00135_),
    .CK(clk),
    .Q(\text_in_r[101] ),
    .QN(_17325_));
 DFF_X1 _34931_ (.D(_00136_),
    .CK(clk),
    .Q(\text_in_r[102] ),
    .QN(_17326_));
 DFF_X1 _34932_ (.D(_00137_),
    .CK(clk),
    .Q(\text_in_r[103] ),
    .QN(_17327_));
 DFF_X1 _34933_ (.D(_00138_),
    .CK(clk),
    .Q(\text_in_r[104] ),
    .QN(_17328_));
 DFF_X1 _34934_ (.D(_00139_),
    .CK(clk),
    .Q(\text_in_r[105] ),
    .QN(_17329_));
 DFF_X1 _34935_ (.D(_00140_),
    .CK(clk),
    .Q(\text_in_r[106] ),
    .QN(_17330_));
 DFF_X1 _34936_ (.D(_00141_),
    .CK(clk),
    .Q(\text_in_r[107] ),
    .QN(_17331_));
 DFF_X1 _34937_ (.D(_00142_),
    .CK(clk),
    .Q(\text_in_r[108] ),
    .QN(_17332_));
 DFF_X1 _34938_ (.D(_00143_),
    .CK(clk),
    .Q(\text_in_r[109] ),
    .QN(_17333_));
 DFF_X1 _34939_ (.D(_00145_),
    .CK(clk),
    .Q(\text_in_r[110] ),
    .QN(_17334_));
 DFF_X1 _34940_ (.D(_00146_),
    .CK(clk),
    .Q(\text_in_r[111] ),
    .QN(_17335_));
 DFF_X1 _34941_ (.D(_00147_),
    .CK(clk),
    .Q(\text_in_r[112] ),
    .QN(_17336_));
 DFF_X1 _34942_ (.D(_00148_),
    .CK(clk),
    .Q(\text_in_r[113] ),
    .QN(_17337_));
 DFF_X1 _34943_ (.D(_00149_),
    .CK(clk),
    .Q(\text_in_r[114] ),
    .QN(_17338_));
 DFF_X1 _34944_ (.D(_00150_),
    .CK(clk),
    .Q(\text_in_r[115] ),
    .QN(_17339_));
 DFF_X1 _34945_ (.D(_00151_),
    .CK(clk),
    .Q(\text_in_r[116] ),
    .QN(_17340_));
 DFF_X1 _34946_ (.D(_00152_),
    .CK(clk),
    .Q(\text_in_r[117] ),
    .QN(_17341_));
 DFF_X1 _34947_ (.D(_00153_),
    .CK(clk),
    .Q(\text_in_r[118] ),
    .QN(_17342_));
 DFF_X1 _34948_ (.D(_00154_),
    .CK(clk),
    .Q(\text_in_r[119] ),
    .QN(_17343_));
 DFF_X1 _34949_ (.D(_00156_),
    .CK(clk),
    .Q(\text_in_r[120] ),
    .QN(_17344_));
 DFF_X1 _34950_ (.D(_00157_),
    .CK(clk),
    .Q(\text_in_r[121] ),
    .QN(_17345_));
 DFF_X1 _34951_ (.D(_00158_),
    .CK(clk),
    .Q(\text_in_r[122] ),
    .QN(_17346_));
 DFF_X1 _34952_ (.D(_00159_),
    .CK(clk),
    .Q(\text_in_r[123] ),
    .QN(_17347_));
 DFF_X1 _34953_ (.D(_00160_),
    .CK(clk),
    .Q(\text_in_r[124] ),
    .QN(_17348_));
 DFF_X1 _34954_ (.D(_00161_),
    .CK(clk),
    .Q(\text_in_r[125] ),
    .QN(_17349_));
 DFF_X1 _34955_ (.D(_00162_),
    .CK(clk),
    .Q(\text_in_r[126] ),
    .QN(_17350_));
 DFF_X1 _34956_ (.D(_00163_),
    .CK(clk),
    .Q(\text_in_r[127] ),
    .QN(_17351_));
 DFF_X1 _34957_ (.D(net2),
    .CK(clk),
    .Q(ld_r),
    .QN(_17352_));
 DFF_X1 _34958_ (.D(_00125_),
    .CK(clk),
    .Q(\sa33[0] ),
    .QN(_17353_));
 DFF_X1 _34959_ (.D(_00126_),
    .CK(clk),
    .Q(\sa33[1] ),
    .QN(_17354_));
 DFF_X1 _34960_ (.D(_00127_),
    .CK(clk),
    .Q(\sa33[2] ),
    .QN(_17355_));
 DFF_X1 _34961_ (.D(_00128_),
    .CK(clk),
    .Q(\sa33[3] ),
    .QN(_17356_));
 DFF_X1 _34962_ (.D(_00129_),
    .CK(clk),
    .Q(\sa33[4] ),
    .QN(_17357_));
 DFF_X1 _34963_ (.D(_00130_),
    .CK(clk),
    .Q(\sa33[5] ),
    .QN(_17358_));
 DFF_X1 _34964_ (.D(_00131_),
    .CK(clk),
    .Q(\sa33[6] ),
    .QN(_17359_));
 DFF_X1 _34965_ (.D(_00132_),
    .CK(clk),
    .Q(\sa33[7] ),
    .QN(_17360_));
 DFF_X1 _34966_ (.D(_00093_),
    .CK(clk),
    .Q(\sa23[0] ),
    .QN(_17361_));
 DFF_X1 _34967_ (.D(_00094_),
    .CK(clk),
    .Q(\sa23[1] ),
    .QN(_17362_));
 DFF_X1 _34968_ (.D(_00095_),
    .CK(clk),
    .Q(\sa23[2] ),
    .QN(_17363_));
 DFF_X1 _34969_ (.D(_00096_),
    .CK(clk),
    .Q(\sa23[3] ),
    .QN(_17364_));
 DFF_X1 _34970_ (.D(_00097_),
    .CK(clk),
    .Q(\sa23[4] ),
    .QN(_17365_));
 DFF_X1 _34971_ (.D(_00098_),
    .CK(clk),
    .Q(\sa23[5] ),
    .QN(_17366_));
 DFF_X1 _34972_ (.D(_00099_),
    .CK(clk),
    .Q(\sa23[6] ),
    .QN(_17367_));
 DFF_X1 _34973_ (.D(_00100_),
    .CK(clk),
    .Q(\sa23[7] ),
    .QN(_17368_));
 DFF_X1 _34974_ (.D(_00061_),
    .CK(clk),
    .Q(\sa13[0] ),
    .QN(_17369_));
 DFF_X1 _34975_ (.D(_00062_),
    .CK(clk),
    .Q(\sa13[1] ),
    .QN(_17370_));
 DFF_X1 _34976_ (.D(_00063_),
    .CK(clk),
    .Q(\sa13[2] ),
    .QN(_17371_));
 DFF_X1 _34977_ (.D(_00064_),
    .CK(clk),
    .Q(\sa13[3] ),
    .QN(_17372_));
 DFF_X1 _34978_ (.D(_00065_),
    .CK(clk),
    .Q(\sa13[4] ),
    .QN(_17373_));
 DFF_X1 _34979_ (.D(_00066_),
    .CK(clk),
    .Q(\sa13[5] ),
    .QN(_17374_));
 DFF_X1 _34980_ (.D(_00067_),
    .CK(clk),
    .Q(\sa13[6] ),
    .QN(_17375_));
 DFF_X1 _34981_ (.D(_00068_),
    .CK(clk),
    .Q(\sa13[7] ),
    .QN(_17376_));
 DFF_X1 _34982_ (.D(_00029_),
    .CK(clk),
    .Q(\sa03[0] ),
    .QN(_17377_));
 DFF_X1 _34983_ (.D(_00030_),
    .CK(clk),
    .Q(\sa03[1] ),
    .QN(_17378_));
 DFF_X1 _34984_ (.D(_00031_),
    .CK(clk),
    .Q(\sa03[2] ),
    .QN(_17379_));
 DFF_X1 _34985_ (.D(_00032_),
    .CK(clk),
    .Q(\sa03[3] ),
    .QN(_17380_));
 DFF_X1 _34986_ (.D(_00033_),
    .CK(clk),
    .Q(\sa03[4] ),
    .QN(_17381_));
 DFF_X1 _34987_ (.D(_00034_),
    .CK(clk),
    .Q(\sa03[5] ),
    .QN(_17382_));
 DFF_X1 _34988_ (.D(_00035_),
    .CK(clk),
    .Q(\sa03[6] ),
    .QN(_17383_));
 DFF_X1 _34989_ (.D(_00036_),
    .CK(clk),
    .Q(\sa03[7] ),
    .QN(_17384_));
 DFF_X1 _34990_ (.D(_00117_),
    .CK(clk),
    .Q(\sa32[0] ),
    .QN(_17385_));
 DFF_X1 _34991_ (.D(_00118_),
    .CK(clk),
    .Q(\sa32[1] ),
    .QN(_17386_));
 DFF_X1 _34992_ (.D(_00119_),
    .CK(clk),
    .Q(\sa32[2] ),
    .QN(_17387_));
 DFF_X1 _34993_ (.D(_00120_),
    .CK(clk),
    .Q(\sa32[3] ),
    .QN(_17388_));
 DFF_X1 _34994_ (.D(_00121_),
    .CK(clk),
    .Q(\sa32[4] ),
    .QN(_17389_));
 DFF_X1 _34995_ (.D(_00122_),
    .CK(clk),
    .Q(\sa32[5] ),
    .QN(_17390_));
 DFF_X1 _34996_ (.D(_00123_),
    .CK(clk),
    .Q(\sa32[6] ),
    .QN(_17391_));
 DFF_X1 _34997_ (.D(_00124_),
    .CK(clk),
    .Q(\sa32[7] ),
    .QN(_17392_));
 DFF_X1 _34998_ (.D(_00085_),
    .CK(clk),
    .Q(\sa22[0] ),
    .QN(_17393_));
 DFF_X1 _34999_ (.D(_00086_),
    .CK(clk),
    .Q(\sa22[1] ),
    .QN(_17394_));
 DFF_X1 _35000_ (.D(_00087_),
    .CK(clk),
    .Q(\sa22[2] ),
    .QN(_17395_));
 DFF_X1 _35001_ (.D(_00088_),
    .CK(clk),
    .Q(\sa22[3] ),
    .QN(_17396_));
 DFF_X1 _35002_ (.D(_00089_),
    .CK(clk),
    .Q(\sa22[4] ),
    .QN(_17397_));
 DFF_X1 _35003_ (.D(_00090_),
    .CK(clk),
    .Q(\sa22[5] ),
    .QN(_17398_));
 DFF_X1 _35004_ (.D(_00091_),
    .CK(clk),
    .Q(\sa22[6] ),
    .QN(_17399_));
 DFF_X1 _35005_ (.D(_00092_),
    .CK(clk),
    .Q(\sa22[7] ),
    .QN(_17400_));
 DFF_X1 _35006_ (.D(_00053_),
    .CK(clk),
    .Q(\sa12[0] ),
    .QN(_17401_));
 DFF_X1 _35007_ (.D(_00054_),
    .CK(clk),
    .Q(\sa12[1] ),
    .QN(_17402_));
 DFF_X1 _35008_ (.D(_00055_),
    .CK(clk),
    .Q(\sa12[2] ),
    .QN(_17403_));
 DFF_X1 _35009_ (.D(_00056_),
    .CK(clk),
    .Q(\sa12[3] ),
    .QN(_17404_));
 DFF_X1 _35010_ (.D(_00057_),
    .CK(clk),
    .Q(\sa12[4] ),
    .QN(_17405_));
 DFF_X1 _35011_ (.D(_00058_),
    .CK(clk),
    .Q(\sa12[5] ),
    .QN(_17406_));
 DFF_X1 _35012_ (.D(_00059_),
    .CK(clk),
    .Q(\sa12[6] ),
    .QN(_17407_));
 DFF_X1 _35013_ (.D(_00060_),
    .CK(clk),
    .Q(\sa12[7] ),
    .QN(_17408_));
 DFF_X1 _35014_ (.D(_00021_),
    .CK(clk),
    .Q(\sa02[0] ),
    .QN(_17409_));
 DFF_X1 _35015_ (.D(_00022_),
    .CK(clk),
    .Q(\sa02[1] ),
    .QN(_17410_));
 DFF_X1 _35016_ (.D(_00023_),
    .CK(clk),
    .Q(\sa02[2] ),
    .QN(_17411_));
 DFF_X1 _35017_ (.D(_00024_),
    .CK(clk),
    .Q(\sa02[3] ),
    .QN(_17412_));
 DFF_X1 _35018_ (.D(_00025_),
    .CK(clk),
    .Q(\sa02[4] ),
    .QN(_17413_));
 DFF_X1 _35019_ (.D(_00026_),
    .CK(clk),
    .Q(\sa02[5] ),
    .QN(_17414_));
 DFF_X1 _35020_ (.D(_00027_),
    .CK(clk),
    .Q(\sa02[6] ),
    .QN(_17415_));
 DFF_X1 _35021_ (.D(_00028_),
    .CK(clk),
    .Q(\sa02[7] ),
    .QN(_17416_));
 DFF_X1 _35022_ (.D(_00109_),
    .CK(clk),
    .Q(\sa31[0] ),
    .QN(_17417_));
 DFF_X1 _35023_ (.D(_00110_),
    .CK(clk),
    .Q(\sa31[1] ),
    .QN(_17418_));
 DFF_X1 _35024_ (.D(_00111_),
    .CK(clk),
    .Q(\sa31[2] ),
    .QN(_17419_));
 DFF_X1 _35025_ (.D(_00112_),
    .CK(clk),
    .Q(\sa31[3] ),
    .QN(_17420_));
 DFF_X1 _35026_ (.D(_00113_),
    .CK(clk),
    .Q(\sa31[4] ),
    .QN(_17421_));
 DFF_X1 _35027_ (.D(_00114_),
    .CK(clk),
    .Q(\sa31[5] ),
    .QN(_17422_));
 DFF_X1 _35028_ (.D(_00115_),
    .CK(clk),
    .Q(\sa31[6] ),
    .QN(_17423_));
 DFF_X1 _35029_ (.D(_00116_),
    .CK(clk),
    .Q(\sa31[7] ),
    .QN(_17424_));
 DFF_X1 _35030_ (.D(_00077_),
    .CK(clk),
    .Q(\sa21[0] ),
    .QN(_17425_));
 DFF_X1 _35031_ (.D(_00078_),
    .CK(clk),
    .Q(\sa21[1] ),
    .QN(_17426_));
 DFF_X1 _35032_ (.D(_00079_),
    .CK(clk),
    .Q(\sa21[2] ),
    .QN(_17427_));
 DFF_X1 _35033_ (.D(_00080_),
    .CK(clk),
    .Q(\sa21[3] ),
    .QN(_17428_));
 DFF_X1 _35034_ (.D(_00081_),
    .CK(clk),
    .Q(\sa21[4] ),
    .QN(_17429_));
 DFF_X1 _35035_ (.D(_00082_),
    .CK(clk),
    .Q(\sa21[5] ),
    .QN(_17430_));
 DFF_X1 _35036_ (.D(_00083_),
    .CK(clk),
    .Q(\sa21[6] ),
    .QN(_17431_));
 DFF_X1 _35037_ (.D(_00084_),
    .CK(clk),
    .Q(\sa21[7] ),
    .QN(_17432_));
 DFF_X1 _35038_ (.D(_00045_),
    .CK(clk),
    .Q(\sa11[0] ),
    .QN(_17433_));
 DFF_X1 _35039_ (.D(_00046_),
    .CK(clk),
    .Q(\sa11[1] ),
    .QN(_17434_));
 DFF_X1 _35040_ (.D(_00047_),
    .CK(clk),
    .Q(\sa11[2] ),
    .QN(_17435_));
 DFF_X1 _35041_ (.D(_00048_),
    .CK(clk),
    .Q(\sa11[3] ),
    .QN(_17436_));
 DFF_X1 _35042_ (.D(_00049_),
    .CK(clk),
    .Q(\sa11[4] ),
    .QN(_17437_));
 DFF_X1 _35043_ (.D(_00050_),
    .CK(clk),
    .Q(\sa11[5] ),
    .QN(_17438_));
 DFF_X1 _35044_ (.D(_00051_),
    .CK(clk),
    .Q(\sa11[6] ),
    .QN(_17439_));
 DFF_X1 _35045_ (.D(_00052_),
    .CK(clk),
    .Q(\sa11[7] ),
    .QN(_17440_));
 DFF_X1 _35046_ (.D(_00013_),
    .CK(clk),
    .Q(\sa01[0] ),
    .QN(_17441_));
 DFF_X1 _35047_ (.D(_00014_),
    .CK(clk),
    .Q(\sa01[1] ),
    .QN(_17442_));
 DFF_X1 _35048_ (.D(_00015_),
    .CK(clk),
    .Q(\sa01[2] ),
    .QN(_17443_));
 DFF_X1 _35049_ (.D(_00016_),
    .CK(clk),
    .Q(\sa01[3] ),
    .QN(_17444_));
 DFF_X1 _35050_ (.D(_00017_),
    .CK(clk),
    .Q(\sa01[4] ),
    .QN(_17445_));
 DFF_X1 _35051_ (.D(_00018_),
    .CK(clk),
    .Q(\sa01[5] ),
    .QN(_17446_));
 DFF_X1 _35052_ (.D(_00019_),
    .CK(clk),
    .Q(\sa01[6] ),
    .QN(_17447_));
 DFF_X1 _35053_ (.D(_00020_),
    .CK(clk),
    .Q(\sa01[7] ),
    .QN(_17448_));
 DFF_X1 _35054_ (.D(_00101_),
    .CK(clk),
    .Q(\sa30[0] ),
    .QN(_17449_));
 DFF_X1 _35055_ (.D(_00102_),
    .CK(clk),
    .Q(\sa30[1] ),
    .QN(_17450_));
 DFF_X1 _35056_ (.D(_00103_),
    .CK(clk),
    .Q(\sa30[2] ),
    .QN(_17451_));
 DFF_X1 _35057_ (.D(_00104_),
    .CK(clk),
    .Q(\sa30[3] ),
    .QN(_17452_));
 DFF_X1 _35058_ (.D(_00105_),
    .CK(clk),
    .Q(\sa30[4] ),
    .QN(_17453_));
 DFF_X1 _35059_ (.D(_00106_),
    .CK(clk),
    .Q(\sa30[5] ),
    .QN(_17454_));
 DFF_X1 _35060_ (.D(_00107_),
    .CK(clk),
    .Q(\sa30[6] ),
    .QN(_17455_));
 DFF_X1 _35061_ (.D(_00108_),
    .CK(clk),
    .Q(\sa30[7] ),
    .QN(_17456_));
 DFF_X1 _35062_ (.D(_00069_),
    .CK(clk),
    .Q(\sa20[0] ),
    .QN(_17457_));
 DFF_X1 _35063_ (.D(_00070_),
    .CK(clk),
    .Q(\sa20[1] ),
    .QN(_17458_));
 DFF_X1 _35064_ (.D(_00071_),
    .CK(clk),
    .Q(\sa20[2] ),
    .QN(_17459_));
 DFF_X1 _35065_ (.D(_00072_),
    .CK(clk),
    .Q(\sa20[3] ),
    .QN(_17460_));
 DFF_X1 _35066_ (.D(_00073_),
    .CK(clk),
    .Q(\sa20[4] ),
    .QN(_17461_));
 DFF_X1 _35067_ (.D(_00074_),
    .CK(clk),
    .Q(\sa20[5] ),
    .QN(_17462_));
 DFF_X1 _35068_ (.D(_00075_),
    .CK(clk),
    .Q(\sa20[6] ),
    .QN(_17463_));
 DFF_X1 _35069_ (.D(_00076_),
    .CK(clk),
    .Q(\sa20[7] ),
    .QN(_17464_));
 DFF_X1 _35070_ (.D(_00037_),
    .CK(clk),
    .Q(\sa10[0] ),
    .QN(_17465_));
 DFF_X1 _35071_ (.D(_00038_),
    .CK(clk),
    .Q(\sa10[1] ),
    .QN(_17466_));
 DFF_X1 _35072_ (.D(_00039_),
    .CK(clk),
    .Q(\sa10[2] ),
    .QN(_17467_));
 DFF_X1 _35073_ (.D(_00040_),
    .CK(clk),
    .Q(\sa10[3] ),
    .QN(_17468_));
 DFF_X1 _35074_ (.D(_00041_),
    .CK(clk),
    .Q(\sa10[4] ),
    .QN(_17469_));
 DFF_X1 _35075_ (.D(_00042_),
    .CK(clk),
    .Q(\sa10[5] ),
    .QN(_17470_));
 DFF_X1 _35076_ (.D(_00043_),
    .CK(clk),
    .Q(\sa10[6] ),
    .QN(_17471_));
 DFF_X1 _35077_ (.D(_00044_),
    .CK(clk),
    .Q(\sa10[7] ),
    .QN(_17472_));
 DFF_X1 _35078_ (.D(_00005_),
    .CK(clk),
    .Q(\sa00[0] ),
    .QN(_17473_));
 DFF_X1 _35079_ (.D(_00006_),
    .CK(clk),
    .Q(\sa00[1] ),
    .QN(_17474_));
 DFF_X1 _35080_ (.D(_00007_),
    .CK(clk),
    .Q(\sa00[2] ),
    .QN(_17475_));
 DFF_X1 _35081_ (.D(_00008_),
    .CK(clk),
    .Q(\sa00[3] ),
    .QN(_17476_));
 DFF_X1 _35082_ (.D(_00009_),
    .CK(clk),
    .Q(\sa00[4] ),
    .QN(_17477_));
 DFF_X1 _35083_ (.D(_00010_),
    .CK(clk),
    .Q(\sa00[5] ),
    .QN(_17478_));
 DFF_X1 _35084_ (.D(_00011_),
    .CK(clk),
    .Q(\sa00[6] ),
    .QN(_17479_));
 DFF_X1 _35085_ (.D(_00012_),
    .CK(clk),
    .Q(\sa00[7] ),
    .QN(_17480_));
 DFF_X1 _35086_ (.D(_00285_),
    .CK(clk),
    .Q(net267),
    .QN(_17481_));
 DFF_X1 _35087_ (.D(_00286_),
    .CK(clk),
    .Q(net266),
    .QN(_17482_));
 DFF_X1 _35088_ (.D(_00287_),
    .CK(clk),
    .Q(net265),
    .QN(_17483_));
 DFF_X1 _35089_ (.D(_00288_),
    .CK(clk),
    .Q(net264),
    .QN(_17484_));
 DFF_X1 _35090_ (.D(_00289_),
    .CK(clk),
    .Q(net263),
    .QN(_17485_));
 DFF_X1 _35091_ (.D(_00290_),
    .CK(clk),
    .Q(net262),
    .QN(_17486_));
 DFF_X1 _35092_ (.D(_00291_),
    .CK(clk),
    .Q(net261),
    .QN(_17487_));
 DFF_X1 _35093_ (.D(_00292_),
    .CK(clk),
    .Q(net260),
    .QN(_17488_));
 DFF_X1 _35094_ (.D(_00381_),
    .CK(clk),
    .Q(net299),
    .QN(_17489_));
 DFF_X1 _35095_ (.D(_00382_),
    .CK(clk),
    .Q(net298),
    .QN(_17490_));
 DFF_X1 _35096_ (.D(_00383_),
    .CK(clk),
    .Q(net297),
    .QN(_17491_));
 DFF_X1 _35097_ (.D(_00384_),
    .CK(clk),
    .Q(net296),
    .QN(_17492_));
 DFF_X1 _35098_ (.D(_00385_),
    .CK(clk),
    .Q(net295),
    .QN(_17493_));
 DFF_X1 _35099_ (.D(_00386_),
    .CK(clk),
    .Q(net294),
    .QN(_17494_));
 DFF_X1 _35100_ (.D(_00387_),
    .CK(clk),
    .Q(net293),
    .QN(_17495_));
 DFF_X1 _35101_ (.D(_00388_),
    .CK(clk),
    .Q(net292),
    .QN(_17496_));
 DFF_X1 _35102_ (.D(_00341_),
    .CK(clk),
    .Q(net331),
    .QN(_17497_));
 DFF_X1 _35103_ (.D(_00342_),
    .CK(clk),
    .Q(net330),
    .QN(_17498_));
 DFF_X1 _35104_ (.D(_00343_),
    .CK(clk),
    .Q(net329),
    .QN(_17499_));
 DFF_X1 _35105_ (.D(_00344_),
    .CK(clk),
    .Q(net328),
    .QN(_17500_));
 DFF_X1 _35106_ (.D(_00345_),
    .CK(clk),
    .Q(net327),
    .QN(_17501_));
 DFF_X1 _35107_ (.D(_00346_),
    .CK(clk),
    .Q(net326),
    .QN(_17502_));
 DFF_X1 _35108_ (.D(_00347_),
    .CK(clk),
    .Q(net325),
    .QN(_17503_));
 DFF_X1 _35109_ (.D(_00348_),
    .CK(clk),
    .Q(net324),
    .QN(_17504_));
 DFF_X1 _35110_ (.D(_00309_),
    .CK(clk),
    .Q(net363),
    .QN(_17505_));
 DFF_X1 _35111_ (.D(_00310_),
    .CK(clk),
    .Q(net362),
    .QN(_17506_));
 DFF_X1 _35112_ (.D(_00311_),
    .CK(clk),
    .Q(net361),
    .QN(_17507_));
 DFF_X1 _35113_ (.D(_00312_),
    .CK(clk),
    .Q(net360),
    .QN(_17508_));
 DFF_X1 _35114_ (.D(_00313_),
    .CK(clk),
    .Q(net359),
    .QN(_17509_));
 DFF_X1 _35115_ (.D(_00314_),
    .CK(clk),
    .Q(net358),
    .QN(_17510_));
 DFF_X1 _35116_ (.D(_00315_),
    .CK(clk),
    .Q(net357),
    .QN(_17511_));
 DFF_X1 _35117_ (.D(_00316_),
    .CK(clk),
    .Q(net356),
    .QN(_17512_));
 DFF_X1 _35118_ (.D(_00277_),
    .CK(clk),
    .Q(net275),
    .QN(_17513_));
 DFF_X1 _35119_ (.D(_00278_),
    .CK(clk),
    .Q(net274),
    .QN(_17514_));
 DFF_X1 _35120_ (.D(_00279_),
    .CK(clk),
    .Q(net273),
    .QN(_17515_));
 DFF_X1 _35121_ (.D(_00280_),
    .CK(clk),
    .Q(net272),
    .QN(_17516_));
 DFF_X1 _35122_ (.D(_00281_),
    .CK(clk),
    .Q(net271),
    .QN(_17517_));
 DFF_X1 _35123_ (.D(_00282_),
    .CK(clk),
    .Q(net270),
    .QN(_17518_));
 DFF_X1 _35124_ (.D(_00283_),
    .CK(clk),
    .Q(net269),
    .QN(_17519_));
 DFF_X1 _35125_ (.D(_00284_),
    .CK(clk),
    .Q(net268),
    .QN(_17520_));
 DFF_X1 _35126_ (.D(_00373_),
    .CK(clk),
    .Q(net307),
    .QN(_17521_));
 DFF_X1 _35127_ (.D(_00374_),
    .CK(clk),
    .Q(net306),
    .QN(_17522_));
 DFF_X1 _35128_ (.D(_00375_),
    .CK(clk),
    .Q(net305),
    .QN(_17523_));
 DFF_X1 _35129_ (.D(_00376_),
    .CK(clk),
    .Q(net304),
    .QN(_17524_));
 DFF_X1 _35130_ (.D(_00377_),
    .CK(clk),
    .Q(net303),
    .QN(_17525_));
 DFF_X1 _35131_ (.D(_00378_),
    .CK(clk),
    .Q(net302),
    .QN(_17526_));
 DFF_X1 _35132_ (.D(_00379_),
    .CK(clk),
    .Q(net301),
    .QN(_17527_));
 DFF_X1 _35133_ (.D(_00380_),
    .CK(clk),
    .Q(net300),
    .QN(_17528_));
 DFF_X1 _35134_ (.D(_00333_),
    .CK(clk),
    .Q(net339),
    .QN(_17529_));
 DFF_X1 _35135_ (.D(_00334_),
    .CK(clk),
    .Q(net338),
    .QN(_17530_));
 DFF_X1 _35136_ (.D(_00335_),
    .CK(clk),
    .Q(net337),
    .QN(_17531_));
 DFF_X1 _35137_ (.D(_00336_),
    .CK(clk),
    .Q(net336),
    .QN(_17532_));
 DFF_X1 _35138_ (.D(_00337_),
    .CK(clk),
    .Q(net335),
    .QN(_17533_));
 DFF_X1 _35139_ (.D(_00338_),
    .CK(clk),
    .Q(net334),
    .QN(_17534_));
 DFF_X1 _35140_ (.D(_00339_),
    .CK(clk),
    .Q(net333),
    .QN(_17535_));
 DFF_X1 _35141_ (.D(_00340_),
    .CK(clk),
    .Q(net332),
    .QN(_17536_));
 DFF_X1 _35142_ (.D(_00301_),
    .CK(clk),
    .Q(net371),
    .QN(_17537_));
 DFF_X1 _35143_ (.D(_00302_),
    .CK(clk),
    .Q(net370),
    .QN(_17538_));
 DFF_X1 _35144_ (.D(_00303_),
    .CK(clk),
    .Q(net369),
    .QN(_17539_));
 DFF_X1 _35145_ (.D(_00304_),
    .CK(clk),
    .Q(net368),
    .QN(_17540_));
 DFF_X1 _35146_ (.D(_00305_),
    .CK(clk),
    .Q(net367),
    .QN(_17541_));
 DFF_X1 _35147_ (.D(_00306_),
    .CK(clk),
    .Q(net366),
    .QN(_17542_));
 DFF_X1 _35148_ (.D(_00307_),
    .CK(clk),
    .Q(net365),
    .QN(_17543_));
 DFF_X1 _35149_ (.D(_00308_),
    .CK(clk),
    .Q(net364),
    .QN(_17544_));
 DFF_X1 _35150_ (.D(_00269_),
    .CK(clk),
    .Q(net283),
    .QN(_17545_));
 DFF_X1 _35151_ (.D(_00270_),
    .CK(clk),
    .Q(net282),
    .QN(_17546_));
 DFF_X1 _35152_ (.D(_00271_),
    .CK(clk),
    .Q(net281),
    .QN(_17547_));
 DFF_X1 _35153_ (.D(_00272_),
    .CK(clk),
    .Q(net280),
    .QN(_17548_));
 DFF_X1 _35154_ (.D(_00273_),
    .CK(clk),
    .Q(net279),
    .QN(_17549_));
 DFF_X1 _35155_ (.D(_00274_),
    .CK(clk),
    .Q(net278),
    .QN(_17550_));
 DFF_X1 _35156_ (.D(_00275_),
    .CK(clk),
    .Q(net277),
    .QN(_17551_));
 DFF_X1 _35157_ (.D(_00276_),
    .CK(clk),
    .Q(net276),
    .QN(_17552_));
 DFF_X1 _35158_ (.D(_00357_),
    .CK(clk),
    .Q(net315),
    .QN(_17553_));
 DFF_X1 _35159_ (.D(_00358_),
    .CK(clk),
    .Q(net314),
    .QN(_17554_));
 DFF_X1 _35160_ (.D(_00359_),
    .CK(clk),
    .Q(net313),
    .QN(_17555_));
 DFF_X1 _35161_ (.D(_00360_),
    .CK(clk),
    .Q(net312),
    .QN(_17556_));
 DFF_X1 _35162_ (.D(_00361_),
    .CK(clk),
    .Q(net311),
    .QN(_17557_));
 DFF_X1 _35163_ (.D(_00362_),
    .CK(clk),
    .Q(net310),
    .QN(_17558_));
 DFF_X1 _35164_ (.D(_00363_),
    .CK(clk),
    .Q(net309),
    .QN(_17559_));
 DFF_X1 _35165_ (.D(_00364_),
    .CK(clk),
    .Q(net308),
    .QN(_17560_));
 DFF_X1 _35166_ (.D(_00325_),
    .CK(clk),
    .Q(net347),
    .QN(_17561_));
 DFF_X1 _35167_ (.D(_00326_),
    .CK(clk),
    .Q(net346),
    .QN(_17562_));
 DFF_X1 _35168_ (.D(_00327_),
    .CK(clk),
    .Q(net345),
    .QN(_17563_));
 DFF_X1 _35169_ (.D(_00328_),
    .CK(clk),
    .Q(net344),
    .QN(_17564_));
 DFF_X1 _35170_ (.D(_00329_),
    .CK(clk),
    .Q(net343),
    .QN(_17565_));
 DFF_X1 _35171_ (.D(_00330_),
    .CK(clk),
    .Q(net342),
    .QN(_17566_));
 DFF_X1 _35172_ (.D(_00331_),
    .CK(clk),
    .Q(net341),
    .QN(_17567_));
 DFF_X1 _35173_ (.D(_00332_),
    .CK(clk),
    .Q(net340),
    .QN(_17568_));
 DFF_X1 _35174_ (.D(_00293_),
    .CK(clk),
    .Q(net379),
    .QN(_17569_));
 DFF_X1 _35175_ (.D(_00294_),
    .CK(clk),
    .Q(net378),
    .QN(_17570_));
 DFF_X1 _35176_ (.D(_00295_),
    .CK(clk),
    .Q(net377),
    .QN(_17571_));
 DFF_X1 _35177_ (.D(_00296_),
    .CK(clk),
    .Q(net376),
    .QN(_17572_));
 DFF_X1 _35178_ (.D(_00297_),
    .CK(clk),
    .Q(net375),
    .QN(_17573_));
 DFF_X1 _35179_ (.D(_00298_),
    .CK(clk),
    .Q(net374),
    .QN(_17574_));
 DFF_X1 _35180_ (.D(_00299_),
    .CK(clk),
    .Q(net373),
    .QN(_17575_));
 DFF_X1 _35181_ (.D(_00300_),
    .CK(clk),
    .Q(net372),
    .QN(_17576_));
 DFF_X1 _35182_ (.D(_00261_),
    .CK(clk),
    .Q(net291),
    .QN(_17577_));
 DFF_X1 _35183_ (.D(_00262_),
    .CK(clk),
    .Q(net290),
    .QN(_17578_));
 DFF_X1 _35184_ (.D(_00263_),
    .CK(clk),
    .Q(net289),
    .QN(_17579_));
 DFF_X1 _35185_ (.D(_00264_),
    .CK(clk),
    .Q(net288),
    .QN(_17580_));
 DFF_X1 _35186_ (.D(_00265_),
    .CK(clk),
    .Q(net287),
    .QN(_17581_));
 DFF_X1 _35187_ (.D(_00266_),
    .CK(clk),
    .Q(net286),
    .QN(_17582_));
 DFF_X1 _35188_ (.D(_00267_),
    .CK(clk),
    .Q(net285),
    .QN(_17583_));
 DFF_X1 _35189_ (.D(_00268_),
    .CK(clk),
    .Q(net284),
    .QN(_17584_));
 DFF_X1 _35190_ (.D(_00349_),
    .CK(clk),
    .Q(net323),
    .QN(_17585_));
 DFF_X1 _35191_ (.D(_00350_),
    .CK(clk),
    .Q(net322),
    .QN(_17586_));
 DFF_X1 _35192_ (.D(_00351_),
    .CK(clk),
    .Q(net321),
    .QN(_17587_));
 DFF_X1 _35193_ (.D(_00352_),
    .CK(clk),
    .Q(net320),
    .QN(_17588_));
 DFF_X1 _35194_ (.D(_00353_),
    .CK(clk),
    .Q(net319),
    .QN(_17589_));
 DFF_X1 _35195_ (.D(_00354_),
    .CK(clk),
    .Q(net318),
    .QN(_17590_));
 DFF_X1 _35196_ (.D(_00355_),
    .CK(clk),
    .Q(net317),
    .QN(_17591_));
 DFF_X1 _35197_ (.D(_00356_),
    .CK(clk),
    .Q(net316),
    .QN(_17592_));
 DFF_X1 _35198_ (.D(_00317_),
    .CK(clk),
    .Q(net355),
    .QN(_17593_));
 DFF_X1 _35199_ (.D(_00318_),
    .CK(clk),
    .Q(net354),
    .QN(_17594_));
 DFF_X1 _35200_ (.D(_00319_),
    .CK(clk),
    .Q(net353),
    .QN(_17595_));
 DFF_X1 _35201_ (.D(_00320_),
    .CK(clk),
    .Q(net352),
    .QN(_17596_));
 DFF_X1 _35202_ (.D(_00321_),
    .CK(clk),
    .Q(net351),
    .QN(_17597_));
 DFF_X1 _35203_ (.D(_00322_),
    .CK(clk),
    .Q(net350),
    .QN(_17598_));
 DFF_X1 _35204_ (.D(_00323_),
    .CK(clk),
    .Q(net349),
    .QN(_17599_));
 DFF_X1 _35205_ (.D(_00324_),
    .CK(clk),
    .Q(net348),
    .QN(_17600_));
 DFF_X1 _35206_ (.D(_00365_),
    .CK(clk),
    .Q(net387),
    .QN(_17601_));
 DFF_X1 _35207_ (.D(_00366_),
    .CK(clk),
    .Q(net386),
    .QN(_17602_));
 DFF_X1 _35208_ (.D(_00367_),
    .CK(clk),
    .Q(net385),
    .QN(_17603_));
 DFF_X1 _35209_ (.D(_00368_),
    .CK(clk),
    .Q(net384),
    .QN(_17604_));
 DFF_X1 _35210_ (.D(_00369_),
    .CK(clk),
    .Q(net383),
    .QN(_17605_));
 DFF_X1 _35211_ (.D(_00370_),
    .CK(clk),
    .Q(net382),
    .QN(_17606_));
 DFF_X1 _35212_ (.D(_00371_),
    .CK(clk),
    .Q(net381),
    .QN(_17607_));
 DFF_X1 _35213_ (.D(_00372_),
    .CK(clk),
    .Q(net380),
    .QN(_17608_));
 DFF_X1 _35214_ (.D(_00459_),
    .CK(clk),
    .Q(\u0.w[0][0] ),
    .QN(_00389_));
 DFF_X1 _35215_ (.D(_00470_),
    .CK(clk),
    .Q(\u0.w[0][1] ),
    .QN(_00390_));
 DFF_X1 _35216_ (.D(_00481_),
    .CK(clk),
    .Q(\u0.w[0][2] ),
    .QN(_00392_));
 DFF_X1 _35217_ (.D(_00484_),
    .CK(clk),
    .Q(\u0.w[0][3] ),
    .QN(_00393_));
 DFF_X1 _35218_ (.D(_00485_),
    .CK(clk),
    .Q(\u0.w[0][4] ),
    .QN(_00394_));
 DFF_X1 _35219_ (.D(_00486_),
    .CK(clk),
    .Q(\u0.w[0][5] ),
    .QN(_00395_));
 DFF_X1 _35220_ (.D(_00487_),
    .CK(clk),
    .Q(\u0.w[0][6] ),
    .QN(_00396_));
 DFF_X1 _35221_ (.D(_00488_),
    .CK(clk),
    .Q(\u0.w[0][7] ),
    .QN(_00397_));
 DFF_X1 _35222_ (.D(_00489_),
    .CK(clk),
    .Q(\u0.w[0][8] ),
    .QN(_00398_));
 DFF_X1 _35223_ (.D(_00490_),
    .CK(clk),
    .Q(\u0.w[0][9] ),
    .QN(_00399_));
 DFF_X1 _35224_ (.D(_00460_),
    .CK(clk),
    .Q(\u0.w[0][10] ),
    .QN(_00400_));
 DFF_X1 _35225_ (.D(_00461_),
    .CK(clk),
    .Q(\u0.w[0][11] ),
    .QN(_00401_));
 DFF_X1 _35226_ (.D(_00462_),
    .CK(clk),
    .Q(\u0.w[0][12] ),
    .QN(_00402_));
 DFF_X1 _35227_ (.D(_00463_),
    .CK(clk),
    .Q(\u0.w[0][13] ),
    .QN(_00403_));
 DFF_X1 _35228_ (.D(_00464_),
    .CK(clk),
    .Q(\u0.w[0][14] ),
    .QN(_00404_));
 DFF_X1 _35229_ (.D(_00465_),
    .CK(clk),
    .Q(\u0.w[0][15] ),
    .QN(_00405_));
 DFF_X1 _35230_ (.D(_00466_),
    .CK(clk),
    .Q(\u0.w[0][16] ),
    .QN(_00406_));
 DFF_X1 _35231_ (.D(_00467_),
    .CK(clk),
    .Q(\u0.w[0][17] ),
    .QN(_00407_));
 DFF_X1 _35232_ (.D(_00468_),
    .CK(clk),
    .Q(\u0.w[0][18] ),
    .QN(_00408_));
 DFF_X1 _35233_ (.D(_00469_),
    .CK(clk),
    .Q(\u0.w[0][19] ),
    .QN(_00409_));
 DFF_X1 _35234_ (.D(_00471_),
    .CK(clk),
    .Q(\u0.w[0][20] ),
    .QN(_00410_));
 DFF_X1 _35235_ (.D(_00472_),
    .CK(clk),
    .Q(\u0.w[0][21] ),
    .QN(_00411_));
 DFF_X1 _35236_ (.D(_00473_),
    .CK(clk),
    .Q(\u0.w[0][22] ),
    .QN(_00412_));
 DFF_X1 _35237_ (.D(_00474_),
    .CK(clk),
    .Q(\u0.w[0][23] ),
    .QN(_00413_));
 DFF_X1 _35238_ (.D(_00475_),
    .CK(clk),
    .Q(\u0.w[0][24] ),
    .QN(_00415_));
 DFF_X1 _35239_ (.D(_00476_),
    .CK(clk),
    .Q(\u0.w[0][25] ),
    .QN(_00417_));
 DFF_X1 _35240_ (.D(_00477_),
    .CK(clk),
    .Q(\u0.w[0][26] ),
    .QN(_00419_));
 DFF_X1 _35241_ (.D(_00478_),
    .CK(clk),
    .Q(\u0.w[0][27] ),
    .QN(_00421_));
 DFF_X1 _35242_ (.D(_00479_),
    .CK(clk),
    .Q(\u0.w[0][28] ),
    .QN(_00423_));
 DFF_X1 _35243_ (.D(_00480_),
    .CK(clk),
    .Q(\u0.w[0][29] ),
    .QN(_00425_));
 DFF_X1 _35244_ (.D(_00482_),
    .CK(clk),
    .Q(\u0.w[0][30] ),
    .QN(_00427_));
 DFF_X1 _35245_ (.D(_00483_),
    .CK(clk),
    .Q(\u0.w[0][31] ),
    .QN(_00429_));
 DFF_X1 _35246_ (.D(_00491_),
    .CK(clk),
    .Q(\u0.w[1][0] ),
    .QN(_17609_));
 DFF_X1 _35247_ (.D(_00502_),
    .CK(clk),
    .Q(\u0.w[1][1] ),
    .QN(_17610_));
 DFF_X1 _35248_ (.D(_00513_),
    .CK(clk),
    .Q(\u0.w[1][2] ),
    .QN(_17611_));
 DFF_X1 _35249_ (.D(_00516_),
    .CK(clk),
    .Q(\u0.w[1][3] ),
    .QN(_17612_));
 DFF_X1 _35250_ (.D(_00517_),
    .CK(clk),
    .Q(\u0.w[1][4] ),
    .QN(_17613_));
 DFF_X1 _35251_ (.D(_00518_),
    .CK(clk),
    .Q(\u0.w[1][5] ),
    .QN(_17614_));
 DFF_X1 _35252_ (.D(_00519_),
    .CK(clk),
    .Q(\u0.w[1][6] ),
    .QN(_17615_));
 DFF_X1 _35253_ (.D(_00520_),
    .CK(clk),
    .Q(\u0.w[1][7] ),
    .QN(_17616_));
 DFF_X1 _35254_ (.D(_00521_),
    .CK(clk),
    .Q(\u0.w[1][8] ),
    .QN(_00438_));
 DFF_X1 _35255_ (.D(_00522_),
    .CK(clk),
    .Q(\u0.w[1][9] ),
    .QN(_17617_));
 DFF_X1 _35256_ (.D(_00492_),
    .CK(clk),
    .Q(\u0.w[1][10] ),
    .QN(_17618_));
 DFF_X1 _35257_ (.D(_00493_),
    .CK(clk),
    .Q(\u0.w[1][11] ),
    .QN(_17619_));
 DFF_X1 _35258_ (.D(_00494_),
    .CK(clk),
    .Q(\u0.w[1][12] ),
    .QN(_17620_));
 DFF_X1 _35259_ (.D(_00495_),
    .CK(clk),
    .Q(\u0.w[1][13] ),
    .QN(_17621_));
 DFF_X1 _35260_ (.D(_00496_),
    .CK(clk),
    .Q(\u0.w[1][14] ),
    .QN(_17622_));
 DFF_X1 _35261_ (.D(_00497_),
    .CK(clk),
    .Q(\u0.w[1][15] ),
    .QN(_17623_));
 DFF_X1 _35262_ (.D(_00498_),
    .CK(clk),
    .Q(\u0.w[1][16] ),
    .QN(_00439_));
 DFF_X1 _35263_ (.D(_00499_),
    .CK(clk),
    .Q(\u0.w[1][17] ),
    .QN(_00440_));
 DFF_X1 _35264_ (.D(_00500_),
    .CK(clk),
    .Q(\u0.w[1][18] ),
    .QN(_17624_));
 DFF_X1 _35265_ (.D(_00501_),
    .CK(clk),
    .Q(\u0.w[1][19] ),
    .QN(_17625_));
 DFF_X1 _35266_ (.D(_00503_),
    .CK(clk),
    .Q(\u0.w[1][20] ),
    .QN(_17626_));
 DFF_X1 _35267_ (.D(_00504_),
    .CK(clk),
    .Q(\u0.w[1][21] ),
    .QN(_00441_));
 DFF_X1 _35268_ (.D(_00505_),
    .CK(clk),
    .Q(\u0.w[1][22] ),
    .QN(_00442_));
 DFF_X1 _35269_ (.D(_00506_),
    .CK(clk),
    .Q(\u0.w[1][23] ),
    .QN(_17627_));
 DFF_X1 _35270_ (.D(_00507_),
    .CK(clk),
    .Q(\u0.w[1][24] ),
    .QN(_00443_));
 DFF_X1 _35271_ (.D(_00508_),
    .CK(clk),
    .Q(\u0.w[1][25] ),
    .QN(_00444_));
 DFF_X1 _35272_ (.D(_00509_),
    .CK(clk),
    .Q(\u0.w[1][26] ),
    .QN(_17628_));
 DFF_X1 _35273_ (.D(_00510_),
    .CK(clk),
    .Q(\u0.w[1][27] ),
    .QN(_17629_));
 DFF_X1 _35274_ (.D(_00511_),
    .CK(clk),
    .Q(\u0.w[1][28] ),
    .QN(_17630_));
 DFF_X1 _35275_ (.D(_00512_),
    .CK(clk),
    .Q(\u0.w[1][29] ),
    .QN(_00445_));
 DFF_X1 _35276_ (.D(_00514_),
    .CK(clk),
    .Q(\u0.w[1][30] ),
    .QN(_00449_));
 DFF_X1 _35277_ (.D(_00515_),
    .CK(clk),
    .Q(\u0.w[1][31] ),
    .QN(_17631_));
 DFF_X1 _35278_ (.D(_00523_),
    .CK(clk),
    .Q(\u0.w[2][0] ),
    .QN(_17632_));
 DFF_X1 _35279_ (.D(_00534_),
    .CK(clk),
    .Q(\u0.w[2][1] ),
    .QN(_17633_));
 DFF_X1 _35280_ (.D(_00545_),
    .CK(clk),
    .Q(\u0.w[2][2] ),
    .QN(_17634_));
 DFF_X1 _35281_ (.D(_00548_),
    .CK(clk),
    .Q(\u0.w[2][3] ),
    .QN(_17635_));
 DFF_X1 _35282_ (.D(_00549_),
    .CK(clk),
    .Q(\u0.w[2][4] ),
    .QN(_17636_));
 DFF_X1 _35283_ (.D(_00550_),
    .CK(clk),
    .Q(\u0.w[2][5] ),
    .QN(_17637_));
 DFF_X1 _35284_ (.D(_00551_),
    .CK(clk),
    .Q(\u0.w[2][6] ),
    .QN(_17638_));
 DFF_X1 _35285_ (.D(_00552_),
    .CK(clk),
    .Q(\u0.w[2][7] ),
    .QN(_17639_));
 DFF_X1 _35286_ (.D(_00553_),
    .CK(clk),
    .Q(\u0.w[2][8] ),
    .QN(_00391_));
 DFF_X1 _35287_ (.D(_00554_),
    .CK(clk),
    .Q(\u0.w[2][9] ),
    .QN(_17640_));
 DFF_X1 _35288_ (.D(_00524_),
    .CK(clk),
    .Q(\u0.w[2][10] ),
    .QN(_17641_));
 DFF_X1 _35289_ (.D(_00525_),
    .CK(clk),
    .Q(\u0.w[2][11] ),
    .QN(_17642_));
 DFF_X1 _35290_ (.D(_00526_),
    .CK(clk),
    .Q(\u0.w[2][12] ),
    .QN(_17643_));
 DFF_X1 _35291_ (.D(_00527_),
    .CK(clk),
    .Q(\u0.w[2][13] ),
    .QN(_17644_));
 DFF_X1 _35292_ (.D(_00528_),
    .CK(clk),
    .Q(\u0.w[2][14] ),
    .QN(_17645_));
 DFF_X1 _35293_ (.D(_00529_),
    .CK(clk),
    .Q(\u0.w[2][15] ),
    .QN(_17646_));
 DFF_X1 _35294_ (.D(_00530_),
    .CK(clk),
    .Q(\u0.w[2][16] ),
    .QN(_00430_));
 DFF_X1 _35295_ (.D(_00531_),
    .CK(clk),
    .Q(\u0.w[2][17] ),
    .QN(_00431_));
 DFF_X1 _35296_ (.D(_00532_),
    .CK(clk),
    .Q(\u0.w[2][18] ),
    .QN(_17647_));
 DFF_X1 _35297_ (.D(_00533_),
    .CK(clk),
    .Q(\u0.w[2][19] ),
    .QN(_17648_));
 DFF_X1 _35298_ (.D(_00535_),
    .CK(clk),
    .Q(\u0.w[2][20] ),
    .QN(_17649_));
 DFF_X1 _35299_ (.D(_00536_),
    .CK(clk),
    .Q(\u0.w[2][21] ),
    .QN(_00432_));
 DFF_X1 _35300_ (.D(_00537_),
    .CK(clk),
    .Q(\u0.w[2][22] ),
    .QN(_00433_));
 DFF_X1 _35301_ (.D(_00538_),
    .CK(clk),
    .Q(\u0.w[2][23] ),
    .QN(_17650_));
 DFF_X1 _35302_ (.D(_00539_),
    .CK(clk),
    .Q(\u0.w[2][24] ),
    .QN(_00434_));
 DFF_X1 _35303_ (.D(_00540_),
    .CK(clk),
    .Q(\u0.w[2][25] ),
    .QN(_00435_));
 DFF_X1 _35304_ (.D(_00541_),
    .CK(clk),
    .Q(\u0.w[2][26] ),
    .QN(_17651_));
 DFF_X1 _35305_ (.D(_00542_),
    .CK(clk),
    .Q(\u0.w[2][27] ),
    .QN(_17652_));
 DFF_X1 _35306_ (.D(_00543_),
    .CK(clk),
    .Q(\u0.w[2][28] ),
    .QN(_17653_));
 DFF_X1 _35307_ (.D(_00544_),
    .CK(clk),
    .Q(\u0.w[2][29] ),
    .QN(_00436_));
 DFF_X1 _35308_ (.D(_00546_),
    .CK(clk),
    .Q(\u0.w[2][30] ),
    .QN(_00437_));
 DFF_X1 _35309_ (.D(_00547_),
    .CK(clk),
    .Q(\u0.w[2][31] ),
    .QN(_17654_));
 BUF_X4 buffer1 (.A(rst),
    .Z(net1));
 BUF_X4 buffer10 (.A(key[120]),
    .Z(net10));
 BUF_X4 buffer100 (.A(key[30]),
    .Z(net100));
 BUF_X4 buffer101 (.A(key[29]),
    .Z(net101));
 BUF_X4 buffer102 (.A(key[28]),
    .Z(net102));
 BUF_X4 buffer103 (.A(key[27]),
    .Z(net103));
 BUF_X4 buffer104 (.A(key[26]),
    .Z(net104));
 BUF_X4 buffer105 (.A(key[25]),
    .Z(net105));
 BUF_X4 buffer106 (.A(key[24]),
    .Z(net106));
 BUF_X4 buffer107 (.A(key[23]),
    .Z(net107));
 BUF_X4 buffer108 (.A(key[22]),
    .Z(net108));
 BUF_X4 buffer109 (.A(key[21]),
    .Z(net109));
 BUF_X4 buffer11 (.A(key[119]),
    .Z(net11));
 BUF_X4 buffer110 (.A(key[20]),
    .Z(net110));
 BUF_X4 buffer111 (.A(key[19]),
    .Z(net111));
 BUF_X4 buffer112 (.A(key[18]),
    .Z(net112));
 BUF_X4 buffer113 (.A(key[17]),
    .Z(net113));
 BUF_X4 buffer114 (.A(key[16]),
    .Z(net114));
 BUF_X4 buffer115 (.A(key[15]),
    .Z(net115));
 BUF_X4 buffer116 (.A(key[14]),
    .Z(net116));
 BUF_X4 buffer117 (.A(key[13]),
    .Z(net117));
 BUF_X4 buffer118 (.A(key[12]),
    .Z(net118));
 BUF_X4 buffer119 (.A(key[11]),
    .Z(net119));
 BUF_X4 buffer12 (.A(key[118]),
    .Z(net12));
 BUF_X4 buffer120 (.A(key[10]),
    .Z(net120));
 BUF_X4 buffer121 (.A(key[9]),
    .Z(net121));
 BUF_X4 buffer122 (.A(key[8]),
    .Z(net122));
 BUF_X4 buffer123 (.A(key[7]),
    .Z(net123));
 BUF_X4 buffer124 (.A(key[6]),
    .Z(net124));
 BUF_X4 buffer125 (.A(key[5]),
    .Z(net125));
 BUF_X4 buffer126 (.A(key[4]),
    .Z(net126));
 BUF_X4 buffer127 (.A(key[3]),
    .Z(net127));
 BUF_X4 buffer128 (.A(key[2]),
    .Z(net128));
 BUF_X4 buffer129 (.A(key[1]),
    .Z(net129));
 BUF_X4 buffer13 (.A(key[117]),
    .Z(net13));
 BUF_X4 buffer130 (.A(key[0]),
    .Z(net130));
 BUF_X4 buffer131 (.A(text_in[127]),
    .Z(net131));
 BUF_X4 buffer132 (.A(text_in[126]),
    .Z(net132));
 BUF_X4 buffer133 (.A(text_in[125]),
    .Z(net133));
 BUF_X4 buffer134 (.A(text_in[124]),
    .Z(net134));
 BUF_X4 buffer135 (.A(text_in[123]),
    .Z(net135));
 BUF_X4 buffer136 (.A(text_in[122]),
    .Z(net136));
 BUF_X4 buffer137 (.A(text_in[121]),
    .Z(net137));
 BUF_X4 buffer138 (.A(text_in[120]),
    .Z(net138));
 BUF_X4 buffer139 (.A(text_in[119]),
    .Z(net139));
 BUF_X4 buffer14 (.A(key[116]),
    .Z(net14));
 BUF_X4 buffer140 (.A(text_in[118]),
    .Z(net140));
 BUF_X4 buffer141 (.A(text_in[117]),
    .Z(net141));
 BUF_X4 buffer142 (.A(text_in[116]),
    .Z(net142));
 BUF_X4 buffer143 (.A(text_in[115]),
    .Z(net143));
 BUF_X4 buffer144 (.A(text_in[114]),
    .Z(net144));
 BUF_X4 buffer145 (.A(text_in[113]),
    .Z(net145));
 BUF_X4 buffer146 (.A(text_in[112]),
    .Z(net146));
 BUF_X4 buffer147 (.A(text_in[111]),
    .Z(net147));
 BUF_X4 buffer148 (.A(text_in[110]),
    .Z(net148));
 BUF_X4 buffer149 (.A(text_in[109]),
    .Z(net149));
 BUF_X4 buffer15 (.A(key[115]),
    .Z(net15));
 BUF_X4 buffer150 (.A(text_in[108]),
    .Z(net150));
 BUF_X4 buffer151 (.A(text_in[107]),
    .Z(net151));
 BUF_X4 buffer152 (.A(text_in[106]),
    .Z(net152));
 BUF_X4 buffer153 (.A(text_in[105]),
    .Z(net153));
 BUF_X4 buffer154 (.A(text_in[104]),
    .Z(net154));
 BUF_X4 buffer155 (.A(text_in[103]),
    .Z(net155));
 BUF_X4 buffer156 (.A(text_in[102]),
    .Z(net156));
 BUF_X4 buffer157 (.A(text_in[101]),
    .Z(net157));
 BUF_X4 buffer158 (.A(text_in[100]),
    .Z(net158));
 BUF_X4 buffer159 (.A(text_in[99]),
    .Z(net159));
 BUF_X4 buffer16 (.A(key[114]),
    .Z(net16));
 BUF_X4 buffer160 (.A(text_in[98]),
    .Z(net160));
 BUF_X4 buffer161 (.A(text_in[97]),
    .Z(net161));
 BUF_X4 buffer162 (.A(text_in[96]),
    .Z(net162));
 BUF_X4 buffer163 (.A(text_in[95]),
    .Z(net163));
 BUF_X4 buffer164 (.A(text_in[94]),
    .Z(net164));
 BUF_X4 buffer165 (.A(text_in[93]),
    .Z(net165));
 BUF_X4 buffer166 (.A(text_in[92]),
    .Z(net166));
 BUF_X4 buffer167 (.A(text_in[91]),
    .Z(net167));
 BUF_X4 buffer168 (.A(text_in[90]),
    .Z(net168));
 BUF_X4 buffer169 (.A(text_in[89]),
    .Z(net169));
 BUF_X4 buffer17 (.A(key[113]),
    .Z(net17));
 BUF_X4 buffer170 (.A(text_in[88]),
    .Z(net170));
 BUF_X4 buffer171 (.A(text_in[87]),
    .Z(net171));
 BUF_X4 buffer172 (.A(text_in[86]),
    .Z(net172));
 BUF_X4 buffer173 (.A(text_in[85]),
    .Z(net173));
 BUF_X4 buffer174 (.A(text_in[84]),
    .Z(net174));
 BUF_X4 buffer175 (.A(text_in[83]),
    .Z(net175));
 BUF_X4 buffer176 (.A(text_in[82]),
    .Z(net176));
 BUF_X4 buffer177 (.A(text_in[81]),
    .Z(net177));
 BUF_X4 buffer178 (.A(text_in[80]),
    .Z(net178));
 BUF_X4 buffer179 (.A(text_in[79]),
    .Z(net179));
 BUF_X4 buffer18 (.A(key[112]),
    .Z(net18));
 BUF_X4 buffer180 (.A(text_in[78]),
    .Z(net180));
 BUF_X4 buffer181 (.A(text_in[77]),
    .Z(net181));
 BUF_X4 buffer182 (.A(text_in[76]),
    .Z(net182));
 BUF_X4 buffer183 (.A(text_in[75]),
    .Z(net183));
 BUF_X4 buffer184 (.A(text_in[74]),
    .Z(net184));
 BUF_X4 buffer185 (.A(text_in[73]),
    .Z(net185));
 BUF_X4 buffer186 (.A(text_in[72]),
    .Z(net186));
 BUF_X4 buffer187 (.A(text_in[71]),
    .Z(net187));
 BUF_X4 buffer188 (.A(text_in[70]),
    .Z(net188));
 BUF_X4 buffer189 (.A(text_in[69]),
    .Z(net189));
 BUF_X4 buffer19 (.A(key[111]),
    .Z(net19));
 BUF_X4 buffer190 (.A(text_in[68]),
    .Z(net190));
 BUF_X4 buffer191 (.A(text_in[67]),
    .Z(net191));
 BUF_X4 buffer192 (.A(text_in[66]),
    .Z(net192));
 BUF_X4 buffer193 (.A(text_in[65]),
    .Z(net193));
 BUF_X4 buffer194 (.A(text_in[64]),
    .Z(net194));
 BUF_X4 buffer195 (.A(text_in[63]),
    .Z(net195));
 BUF_X4 buffer196 (.A(text_in[62]),
    .Z(net196));
 BUF_X4 buffer197 (.A(text_in[61]),
    .Z(net197));
 BUF_X4 buffer198 (.A(text_in[60]),
    .Z(net198));
 BUF_X4 buffer199 (.A(text_in[59]),
    .Z(net199));
 BUF_X4 buffer2 (.A(ld),
    .Z(net2));
 BUF_X4 buffer20 (.A(key[110]),
    .Z(net20));
 BUF_X4 buffer200 (.A(text_in[58]),
    .Z(net200));
 BUF_X4 buffer201 (.A(text_in[57]),
    .Z(net201));
 BUF_X4 buffer202 (.A(text_in[56]),
    .Z(net202));
 BUF_X4 buffer203 (.A(text_in[55]),
    .Z(net203));
 BUF_X4 buffer204 (.A(text_in[54]),
    .Z(net204));
 BUF_X4 buffer205 (.A(text_in[53]),
    .Z(net205));
 BUF_X4 buffer206 (.A(text_in[52]),
    .Z(net206));
 BUF_X4 buffer207 (.A(text_in[51]),
    .Z(net207));
 BUF_X4 buffer208 (.A(text_in[50]),
    .Z(net208));
 BUF_X4 buffer209 (.A(text_in[49]),
    .Z(net209));
 BUF_X4 buffer21 (.A(key[109]),
    .Z(net21));
 BUF_X4 buffer210 (.A(text_in[48]),
    .Z(net210));
 BUF_X4 buffer211 (.A(text_in[47]),
    .Z(net211));
 BUF_X4 buffer212 (.A(text_in[46]),
    .Z(net212));
 BUF_X4 buffer213 (.A(text_in[45]),
    .Z(net213));
 BUF_X4 buffer214 (.A(text_in[44]),
    .Z(net214));
 BUF_X4 buffer215 (.A(text_in[43]),
    .Z(net215));
 BUF_X4 buffer216 (.A(text_in[42]),
    .Z(net216));
 BUF_X4 buffer217 (.A(text_in[41]),
    .Z(net217));
 BUF_X4 buffer218 (.A(text_in[40]),
    .Z(net218));
 BUF_X4 buffer219 (.A(text_in[39]),
    .Z(net219));
 BUF_X4 buffer22 (.A(key[108]),
    .Z(net22));
 BUF_X4 buffer220 (.A(text_in[38]),
    .Z(net220));
 BUF_X4 buffer221 (.A(text_in[37]),
    .Z(net221));
 BUF_X4 buffer222 (.A(text_in[36]),
    .Z(net222));
 BUF_X4 buffer223 (.A(text_in[35]),
    .Z(net223));
 BUF_X4 buffer224 (.A(text_in[34]),
    .Z(net224));
 BUF_X4 buffer225 (.A(text_in[33]),
    .Z(net225));
 BUF_X4 buffer226 (.A(text_in[32]),
    .Z(net226));
 BUF_X4 buffer227 (.A(text_in[31]),
    .Z(net227));
 BUF_X4 buffer228 (.A(text_in[30]),
    .Z(net228));
 BUF_X4 buffer229 (.A(text_in[29]),
    .Z(net229));
 BUF_X4 buffer23 (.A(key[107]),
    .Z(net23));
 BUF_X4 buffer230 (.A(text_in[28]),
    .Z(net230));
 BUF_X4 buffer231 (.A(text_in[27]),
    .Z(net231));
 BUF_X4 buffer232 (.A(text_in[26]),
    .Z(net232));
 BUF_X4 buffer233 (.A(text_in[25]),
    .Z(net233));
 BUF_X4 buffer234 (.A(text_in[24]),
    .Z(net234));
 BUF_X4 buffer235 (.A(text_in[23]),
    .Z(net235));
 BUF_X4 buffer236 (.A(text_in[22]),
    .Z(net236));
 BUF_X4 buffer237 (.A(text_in[21]),
    .Z(net237));
 BUF_X4 buffer238 (.A(text_in[20]),
    .Z(net238));
 BUF_X4 buffer239 (.A(text_in[19]),
    .Z(net239));
 BUF_X4 buffer24 (.A(key[106]),
    .Z(net24));
 BUF_X4 buffer240 (.A(text_in[18]),
    .Z(net240));
 BUF_X4 buffer241 (.A(text_in[17]),
    .Z(net241));
 BUF_X4 buffer242 (.A(text_in[16]),
    .Z(net242));
 BUF_X4 buffer243 (.A(text_in[15]),
    .Z(net243));
 BUF_X4 buffer244 (.A(text_in[14]),
    .Z(net244));
 BUF_X4 buffer245 (.A(text_in[13]),
    .Z(net245));
 BUF_X4 buffer246 (.A(text_in[12]),
    .Z(net246));
 BUF_X4 buffer247 (.A(text_in[11]),
    .Z(net247));
 BUF_X4 buffer248 (.A(text_in[10]),
    .Z(net248));
 BUF_X4 buffer249 (.A(text_in[9]),
    .Z(net249));
 BUF_X4 buffer25 (.A(key[105]),
    .Z(net25));
 BUF_X4 buffer250 (.A(text_in[8]),
    .Z(net250));
 BUF_X4 buffer251 (.A(text_in[7]),
    .Z(net251));
 BUF_X4 buffer252 (.A(text_in[6]),
    .Z(net252));
 BUF_X4 buffer253 (.A(text_in[5]),
    .Z(net253));
 BUF_X4 buffer254 (.A(text_in[4]),
    .Z(net254));
 BUF_X4 buffer255 (.A(text_in[3]),
    .Z(net255));
 BUF_X4 buffer256 (.A(text_in[2]),
    .Z(net256));
 BUF_X4 buffer257 (.A(text_in[1]),
    .Z(net257));
 BUF_X4 buffer258 (.A(text_in[0]),
    .Z(net258));
 BUF_X4 buffer259 (.A(net259),
    .Z(done));
 BUF_X4 buffer26 (.A(key[104]),
    .Z(net26));
 BUF_X4 buffer260 (.A(net260),
    .Z(text_out[127]));
 BUF_X4 buffer261 (.A(net261),
    .Z(text_out[126]));
 BUF_X4 buffer262 (.A(net262),
    .Z(text_out[125]));
 BUF_X4 buffer263 (.A(net263),
    .Z(text_out[124]));
 BUF_X4 buffer264 (.A(net264),
    .Z(text_out[123]));
 BUF_X4 buffer265 (.A(net265),
    .Z(text_out[122]));
 BUF_X4 buffer266 (.A(net266),
    .Z(text_out[121]));
 BUF_X4 buffer267 (.A(net267),
    .Z(text_out[120]));
 BUF_X4 buffer268 (.A(net268),
    .Z(text_out[119]));
 BUF_X4 buffer269 (.A(net269),
    .Z(text_out[118]));
 BUF_X4 buffer27 (.A(key[103]),
    .Z(net27));
 BUF_X4 buffer270 (.A(net270),
    .Z(text_out[117]));
 BUF_X4 buffer271 (.A(net271),
    .Z(text_out[116]));
 BUF_X4 buffer272 (.A(net272),
    .Z(text_out[115]));
 BUF_X4 buffer273 (.A(net273),
    .Z(text_out[114]));
 BUF_X4 buffer274 (.A(net274),
    .Z(text_out[113]));
 BUF_X4 buffer275 (.A(net275),
    .Z(text_out[112]));
 BUF_X4 buffer276 (.A(net276),
    .Z(text_out[111]));
 BUF_X4 buffer277 (.A(net277),
    .Z(text_out[110]));
 BUF_X4 buffer278 (.A(net278),
    .Z(text_out[109]));
 BUF_X4 buffer279 (.A(net279),
    .Z(text_out[108]));
 BUF_X4 buffer28 (.A(key[102]),
    .Z(net28));
 BUF_X4 buffer280 (.A(net280),
    .Z(text_out[107]));
 BUF_X4 buffer281 (.A(net281),
    .Z(text_out[106]));
 BUF_X4 buffer282 (.A(net282),
    .Z(text_out[105]));
 BUF_X4 buffer283 (.A(net283),
    .Z(text_out[104]));
 BUF_X4 buffer284 (.A(net284),
    .Z(text_out[103]));
 BUF_X4 buffer285 (.A(net285),
    .Z(text_out[102]));
 BUF_X4 buffer286 (.A(net286),
    .Z(text_out[101]));
 BUF_X4 buffer287 (.A(net287),
    .Z(text_out[100]));
 BUF_X4 buffer288 (.A(net288),
    .Z(text_out[99]));
 BUF_X4 buffer289 (.A(net289),
    .Z(text_out[98]));
 BUF_X4 buffer29 (.A(key[101]),
    .Z(net29));
 BUF_X4 buffer290 (.A(net290),
    .Z(text_out[97]));
 BUF_X4 buffer291 (.A(net291),
    .Z(text_out[96]));
 BUF_X4 buffer292 (.A(net292),
    .Z(text_out[95]));
 BUF_X4 buffer293 (.A(net293),
    .Z(text_out[94]));
 BUF_X4 buffer294 (.A(net294),
    .Z(text_out[93]));
 BUF_X4 buffer295 (.A(net295),
    .Z(text_out[92]));
 BUF_X4 buffer296 (.A(net296),
    .Z(text_out[91]));
 BUF_X4 buffer297 (.A(net297),
    .Z(text_out[90]));
 BUF_X4 buffer298 (.A(net298),
    .Z(text_out[89]));
 BUF_X4 buffer299 (.A(net299),
    .Z(text_out[88]));
 BUF_X4 buffer3 (.A(key[127]),
    .Z(net3));
 BUF_X4 buffer30 (.A(key[100]),
    .Z(net30));
 BUF_X4 buffer300 (.A(net300),
    .Z(text_out[87]));
 BUF_X4 buffer301 (.A(net301),
    .Z(text_out[86]));
 BUF_X4 buffer302 (.A(net302),
    .Z(text_out[85]));
 BUF_X4 buffer303 (.A(net303),
    .Z(text_out[84]));
 BUF_X4 buffer304 (.A(net304),
    .Z(text_out[83]));
 BUF_X4 buffer305 (.A(net305),
    .Z(text_out[82]));
 BUF_X4 buffer306 (.A(net306),
    .Z(text_out[81]));
 BUF_X4 buffer307 (.A(net307),
    .Z(text_out[80]));
 BUF_X4 buffer308 (.A(net308),
    .Z(text_out[79]));
 BUF_X4 buffer309 (.A(net309),
    .Z(text_out[78]));
 BUF_X4 buffer31 (.A(key[99]),
    .Z(net31));
 BUF_X4 buffer310 (.A(net310),
    .Z(text_out[77]));
 BUF_X4 buffer311 (.A(net311),
    .Z(text_out[76]));
 BUF_X4 buffer312 (.A(net312),
    .Z(text_out[75]));
 BUF_X4 buffer313 (.A(net313),
    .Z(text_out[74]));
 BUF_X4 buffer314 (.A(net314),
    .Z(text_out[73]));
 BUF_X4 buffer315 (.A(net315),
    .Z(text_out[72]));
 BUF_X4 buffer316 (.A(net316),
    .Z(text_out[71]));
 BUF_X4 buffer317 (.A(net317),
    .Z(text_out[70]));
 BUF_X4 buffer318 (.A(net318),
    .Z(text_out[69]));
 BUF_X4 buffer319 (.A(net319),
    .Z(text_out[68]));
 BUF_X4 buffer32 (.A(key[98]),
    .Z(net32));
 BUF_X4 buffer320 (.A(net320),
    .Z(text_out[67]));
 BUF_X4 buffer321 (.A(net321),
    .Z(text_out[66]));
 BUF_X4 buffer322 (.A(net322),
    .Z(text_out[65]));
 BUF_X4 buffer323 (.A(net323),
    .Z(text_out[64]));
 BUF_X4 buffer324 (.A(net324),
    .Z(text_out[63]));
 BUF_X4 buffer325 (.A(net325),
    .Z(text_out[62]));
 BUF_X4 buffer326 (.A(net326),
    .Z(text_out[61]));
 BUF_X4 buffer327 (.A(net327),
    .Z(text_out[60]));
 BUF_X4 buffer328 (.A(net328),
    .Z(text_out[59]));
 BUF_X4 buffer329 (.A(net329),
    .Z(text_out[58]));
 BUF_X4 buffer33 (.A(key[97]),
    .Z(net33));
 BUF_X4 buffer330 (.A(net330),
    .Z(text_out[57]));
 BUF_X4 buffer331 (.A(net331),
    .Z(text_out[56]));
 BUF_X4 buffer332 (.A(net332),
    .Z(text_out[55]));
 BUF_X4 buffer333 (.A(net333),
    .Z(text_out[54]));
 BUF_X4 buffer334 (.A(net334),
    .Z(text_out[53]));
 BUF_X4 buffer335 (.A(net335),
    .Z(text_out[52]));
 BUF_X4 buffer336 (.A(net336),
    .Z(text_out[51]));
 BUF_X4 buffer337 (.A(net337),
    .Z(text_out[50]));
 BUF_X4 buffer338 (.A(net338),
    .Z(text_out[49]));
 BUF_X4 buffer339 (.A(net339),
    .Z(text_out[48]));
 BUF_X4 buffer34 (.A(key[96]),
    .Z(net34));
 BUF_X4 buffer340 (.A(net340),
    .Z(text_out[47]));
 BUF_X4 buffer341 (.A(net341),
    .Z(text_out[46]));
 BUF_X4 buffer342 (.A(net342),
    .Z(text_out[45]));
 BUF_X4 buffer343 (.A(net343),
    .Z(text_out[44]));
 BUF_X4 buffer344 (.A(net344),
    .Z(text_out[43]));
 BUF_X4 buffer345 (.A(net345),
    .Z(text_out[42]));
 BUF_X4 buffer346 (.A(net346),
    .Z(text_out[41]));
 BUF_X4 buffer347 (.A(net347),
    .Z(text_out[40]));
 BUF_X4 buffer348 (.A(net348),
    .Z(text_out[39]));
 BUF_X4 buffer349 (.A(net349),
    .Z(text_out[38]));
 BUF_X4 buffer35 (.A(key[95]),
    .Z(net35));
 BUF_X4 buffer350 (.A(net350),
    .Z(text_out[37]));
 BUF_X4 buffer351 (.A(net351),
    .Z(text_out[36]));
 BUF_X4 buffer352 (.A(net352),
    .Z(text_out[35]));
 BUF_X4 buffer353 (.A(net353),
    .Z(text_out[34]));
 BUF_X4 buffer354 (.A(net354),
    .Z(text_out[33]));
 BUF_X4 buffer355 (.A(net355),
    .Z(text_out[32]));
 BUF_X4 buffer356 (.A(net356),
    .Z(text_out[31]));
 BUF_X4 buffer357 (.A(net357),
    .Z(text_out[30]));
 BUF_X4 buffer358 (.A(net358),
    .Z(text_out[29]));
 BUF_X4 buffer359 (.A(net359),
    .Z(text_out[28]));
 BUF_X4 buffer36 (.A(key[94]),
    .Z(net36));
 BUF_X4 buffer360 (.A(net360),
    .Z(text_out[27]));
 BUF_X4 buffer361 (.A(net361),
    .Z(text_out[26]));
 BUF_X4 buffer362 (.A(net362),
    .Z(text_out[25]));
 BUF_X4 buffer363 (.A(net363),
    .Z(text_out[24]));
 BUF_X4 buffer364 (.A(net364),
    .Z(text_out[23]));
 BUF_X4 buffer365 (.A(net365),
    .Z(text_out[22]));
 BUF_X4 buffer366 (.A(net366),
    .Z(text_out[21]));
 BUF_X4 buffer367 (.A(net367),
    .Z(text_out[20]));
 BUF_X4 buffer368 (.A(net368),
    .Z(text_out[19]));
 BUF_X4 buffer369 (.A(net369),
    .Z(text_out[18]));
 BUF_X4 buffer37 (.A(key[93]),
    .Z(net37));
 BUF_X4 buffer370 (.A(net370),
    .Z(text_out[17]));
 BUF_X4 buffer371 (.A(net371),
    .Z(text_out[16]));
 BUF_X4 buffer372 (.A(net372),
    .Z(text_out[15]));
 BUF_X4 buffer373 (.A(net373),
    .Z(text_out[14]));
 BUF_X4 buffer374 (.A(net374),
    .Z(text_out[13]));
 BUF_X4 buffer375 (.A(net375),
    .Z(text_out[12]));
 BUF_X4 buffer376 (.A(net376),
    .Z(text_out[11]));
 BUF_X4 buffer377 (.A(net377),
    .Z(text_out[10]));
 BUF_X4 buffer378 (.A(net378),
    .Z(text_out[9]));
 BUF_X4 buffer379 (.A(net379),
    .Z(text_out[8]));
 BUF_X4 buffer38 (.A(key[92]),
    .Z(net38));
 BUF_X4 buffer380 (.A(net380),
    .Z(text_out[7]));
 BUF_X4 buffer381 (.A(net381),
    .Z(text_out[6]));
 BUF_X4 buffer382 (.A(net382),
    .Z(text_out[5]));
 BUF_X4 buffer383 (.A(net383),
    .Z(text_out[4]));
 BUF_X4 buffer384 (.A(net384),
    .Z(text_out[3]));
 BUF_X4 buffer385 (.A(net385),
    .Z(text_out[2]));
 BUF_X4 buffer386 (.A(net386),
    .Z(text_out[1]));
 BUF_X4 buffer387 (.A(net387),
    .Z(text_out[0]));
 BUF_X4 buffer39 (.A(key[91]),
    .Z(net39));
 BUF_X4 buffer4 (.A(key[126]),
    .Z(net4));
 BUF_X4 buffer40 (.A(key[90]),
    .Z(net40));
 BUF_X4 buffer41 (.A(key[89]),
    .Z(net41));
 BUF_X4 buffer42 (.A(key[88]),
    .Z(net42));
 BUF_X4 buffer43 (.A(key[87]),
    .Z(net43));
 BUF_X4 buffer44 (.A(key[86]),
    .Z(net44));
 BUF_X4 buffer45 (.A(key[85]),
    .Z(net45));
 BUF_X4 buffer46 (.A(key[84]),
    .Z(net46));
 BUF_X4 buffer47 (.A(key[83]),
    .Z(net47));
 BUF_X4 buffer48 (.A(key[82]),
    .Z(net48));
 BUF_X4 buffer49 (.A(key[81]),
    .Z(net49));
 BUF_X4 buffer5 (.A(key[125]),
    .Z(net5));
 BUF_X4 buffer50 (.A(key[80]),
    .Z(net50));
 BUF_X4 buffer51 (.A(key[79]),
    .Z(net51));
 BUF_X4 buffer52 (.A(key[78]),
    .Z(net52));
 BUF_X4 buffer53 (.A(key[77]),
    .Z(net53));
 BUF_X4 buffer54 (.A(key[76]),
    .Z(net54));
 BUF_X4 buffer55 (.A(key[75]),
    .Z(net55));
 BUF_X4 buffer56 (.A(key[74]),
    .Z(net56));
 BUF_X4 buffer57 (.A(key[73]),
    .Z(net57));
 BUF_X4 buffer58 (.A(key[72]),
    .Z(net58));
 BUF_X4 buffer59 (.A(key[71]),
    .Z(net59));
 BUF_X4 buffer6 (.A(key[124]),
    .Z(net6));
 BUF_X4 buffer60 (.A(key[70]),
    .Z(net60));
 BUF_X4 buffer61 (.A(key[69]),
    .Z(net61));
 BUF_X4 buffer62 (.A(key[68]),
    .Z(net62));
 BUF_X4 buffer63 (.A(key[67]),
    .Z(net63));
 BUF_X4 buffer64 (.A(key[66]),
    .Z(net64));
 BUF_X4 buffer65 (.A(key[65]),
    .Z(net65));
 BUF_X4 buffer66 (.A(key[64]),
    .Z(net66));
 BUF_X4 buffer67 (.A(key[63]),
    .Z(net67));
 BUF_X4 buffer68 (.A(key[62]),
    .Z(net68));
 BUF_X4 buffer69 (.A(key[61]),
    .Z(net69));
 BUF_X4 buffer7 (.A(key[123]),
    .Z(net7));
 BUF_X4 buffer70 (.A(key[60]),
    .Z(net70));
 BUF_X4 buffer71 (.A(key[59]),
    .Z(net71));
 BUF_X4 buffer72 (.A(key[58]),
    .Z(net72));
 BUF_X4 buffer73 (.A(key[57]),
    .Z(net73));
 BUF_X4 buffer74 (.A(key[56]),
    .Z(net74));
 BUF_X4 buffer75 (.A(key[55]),
    .Z(net75));
 BUF_X4 buffer76 (.A(key[54]),
    .Z(net76));
 BUF_X4 buffer77 (.A(key[53]),
    .Z(net77));
 BUF_X4 buffer78 (.A(key[52]),
    .Z(net78));
 BUF_X4 buffer79 (.A(key[51]),
    .Z(net79));
 BUF_X4 buffer8 (.A(key[122]),
    .Z(net8));
 BUF_X4 buffer80 (.A(key[50]),
    .Z(net80));
 BUF_X4 buffer81 (.A(key[49]),
    .Z(net81));
 BUF_X4 buffer82 (.A(key[48]),
    .Z(net82));
 BUF_X4 buffer83 (.A(key[47]),
    .Z(net83));
 BUF_X4 buffer84 (.A(key[46]),
    .Z(net84));
 BUF_X4 buffer85 (.A(key[45]),
    .Z(net85));
 BUF_X4 buffer86 (.A(key[44]),
    .Z(net86));
 BUF_X4 buffer87 (.A(key[43]),
    .Z(net87));
 BUF_X4 buffer88 (.A(key[42]),
    .Z(net88));
 BUF_X4 buffer89 (.A(key[41]),
    .Z(net89));
 BUF_X4 buffer9 (.A(key[121]),
    .Z(net9));
 BUF_X4 buffer90 (.A(key[40]),
    .Z(net90));
 BUF_X4 buffer91 (.A(key[39]),
    .Z(net91));
 BUF_X4 buffer92 (.A(key[38]),
    .Z(net92));
 BUF_X4 buffer93 (.A(key[37]),
    .Z(net93));
 BUF_X4 buffer94 (.A(key[36]),
    .Z(net94));
 BUF_X4 buffer95 (.A(key[35]),
    .Z(net95));
 BUF_X4 buffer96 (.A(key[34]),
    .Z(net96));
 BUF_X4 buffer97 (.A(key[33]),
    .Z(net97));
 BUF_X4 buffer98 (.A(key[32]),
    .Z(net98));
 BUF_X4 buffer99 (.A(key[31]),
    .Z(net99));
endmodule
