VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_64x32
  FOREIGN fakeram45_64x32 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 19.190 BY 56.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.785 0.070 1.855 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.205 0.070 2.275 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.625 0.070 2.695 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.045 0.070 3.115 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.465 0.070 3.535 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.885 0.070 3.955 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.305 0.070 4.375 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.725 0.070 4.795 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.145 0.070 5.215 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.565 0.070 5.635 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.985 0.070 6.055 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.405 0.070 6.475 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.825 0.070 6.895 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.245 0.070 7.315 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.665 0.070 7.735 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.085 0.070 8.155 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.505 0.070 8.575 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.925 0.070 8.995 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.345 0.070 9.415 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.765 0.070 9.835 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.185 0.070 10.255 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.605 0.070 10.675 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.025 0.070 11.095 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.445 0.070 11.515 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.865 0.070 11.935 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.285 0.070 12.355 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.705 0.070 12.775 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.125 0.070 13.195 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.545 0.070 13.615 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.965 0.070 14.035 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.385 0.070 14.455 ;
    END
  END w_mask_in[31]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.625 0.070 16.695 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.045 0.070 17.115 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.465 0.070 17.535 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.885 0.070 17.955 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.305 0.070 18.375 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.725 0.070 18.795 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.145 0.070 19.215 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.565 0.070 19.635 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.985 0.070 20.055 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.405 0.070 20.475 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.825 0.070 20.895 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.245 0.070 21.315 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.665 0.070 21.735 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.085 0.070 22.155 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.505 0.070 22.575 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.925 0.070 22.995 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.345 0.070 23.415 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.765 0.070 23.835 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.185 0.070 24.255 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.605 0.070 24.675 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.025 0.070 25.095 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.445 0.070 25.515 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.865 0.070 25.935 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.285 0.070 26.355 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.705 0.070 26.775 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.125 0.070 27.195 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.545 0.070 27.615 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.965 0.070 28.035 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.385 0.070 28.455 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.805 0.070 28.875 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.225 0.070 29.295 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.645 0.070 29.715 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.885 0.070 31.955 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.305 0.070 32.375 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.725 0.070 32.795 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.145 0.070 33.215 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.565 0.070 33.635 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.985 0.070 34.055 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.405 0.070 34.475 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.825 0.070 34.895 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.245 0.070 35.315 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.665 0.070 35.735 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.085 0.070 36.155 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.505 0.070 36.575 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.925 0.070 36.995 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.185 0.070 38.255 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.025 0.070 39.095 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.705 0.070 40.775 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.545 0.070 41.615 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.385 0.070 42.455 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.805 0.070 42.875 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.065 0.070 44.135 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.905 0.070 44.975 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.145 0.070 47.215 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.565 0.070 47.635 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.985 0.070 48.055 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.405 0.070 48.475 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.825 0.070 48.895 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.245 0.070 49.315 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.485 0.070 51.555 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.905 0.070 51.975 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.325 0.070 52.395 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 54.600 ;
      RECT 3.500 1.400 3.780 54.600 ;
      RECT 5.740 1.400 6.020 54.600 ;
      RECT 7.980 1.400 8.260 54.600 ;
      RECT 10.220 1.400 10.500 54.600 ;
      RECT 12.460 1.400 12.740 54.600 ;
      RECT 14.700 1.400 14.980 54.600 ;
      RECT 16.940 1.400 17.220 54.600 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 54.600 ;
      RECT 4.620 1.400 4.900 54.600 ;
      RECT 6.860 1.400 7.140 54.600 ;
      RECT 9.100 1.400 9.380 54.600 ;
      RECT 11.340 1.400 11.620 54.600 ;
      RECT 13.580 1.400 13.860 54.600 ;
      RECT 15.820 1.400 16.100 54.600 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 19.190 56.000 ;
    LAYER metal2 ;
    RECT 0 0 19.190 56.000 ;
    LAYER metal3 ;
    RECT 0.070 0 19.190 56.000 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 1.785 ;
    RECT 0 1.855 0.070 2.205 ;
    RECT 0 2.275 0.070 2.625 ;
    RECT 0 2.695 0.070 3.045 ;
    RECT 0 3.115 0.070 3.465 ;
    RECT 0 3.535 0.070 3.885 ;
    RECT 0 3.955 0.070 4.305 ;
    RECT 0 4.375 0.070 4.725 ;
    RECT 0 4.795 0.070 5.145 ;
    RECT 0 5.215 0.070 5.565 ;
    RECT 0 5.635 0.070 5.985 ;
    RECT 0 6.055 0.070 6.405 ;
    RECT 0 6.475 0.070 6.825 ;
    RECT 0 6.895 0.070 7.245 ;
    RECT 0 7.315 0.070 7.665 ;
    RECT 0 7.735 0.070 8.085 ;
    RECT 0 8.155 0.070 8.505 ;
    RECT 0 8.575 0.070 8.925 ;
    RECT 0 8.995 0.070 9.345 ;
    RECT 0 9.415 0.070 9.765 ;
    RECT 0 9.835 0.070 10.185 ;
    RECT 0 10.255 0.070 10.605 ;
    RECT 0 10.675 0.070 11.025 ;
    RECT 0 11.095 0.070 11.445 ;
    RECT 0 11.515 0.070 11.865 ;
    RECT 0 11.935 0.070 12.285 ;
    RECT 0 12.355 0.070 12.705 ;
    RECT 0 12.775 0.070 13.125 ;
    RECT 0 13.195 0.070 13.545 ;
    RECT 0 13.615 0.070 13.965 ;
    RECT 0 14.035 0.070 14.385 ;
    RECT 0 14.455 0.070 16.625 ;
    RECT 0 16.695 0.070 17.045 ;
    RECT 0 17.115 0.070 17.465 ;
    RECT 0 17.535 0.070 17.885 ;
    RECT 0 17.955 0.070 18.305 ;
    RECT 0 18.375 0.070 18.725 ;
    RECT 0 18.795 0.070 19.145 ;
    RECT 0 19.215 0.070 19.565 ;
    RECT 0 19.635 0.070 19.985 ;
    RECT 0 20.055 0.070 20.405 ;
    RECT 0 20.475 0.070 20.825 ;
    RECT 0 20.895 0.070 21.245 ;
    RECT 0 21.315 0.070 21.665 ;
    RECT 0 21.735 0.070 22.085 ;
    RECT 0 22.155 0.070 22.505 ;
    RECT 0 22.575 0.070 22.925 ;
    RECT 0 22.995 0.070 23.345 ;
    RECT 0 23.415 0.070 23.765 ;
    RECT 0 23.835 0.070 24.185 ;
    RECT 0 24.255 0.070 24.605 ;
    RECT 0 24.675 0.070 25.025 ;
    RECT 0 25.095 0.070 25.445 ;
    RECT 0 25.515 0.070 25.865 ;
    RECT 0 25.935 0.070 26.285 ;
    RECT 0 26.355 0.070 26.705 ;
    RECT 0 26.775 0.070 27.125 ;
    RECT 0 27.195 0.070 27.545 ;
    RECT 0 27.615 0.070 27.965 ;
    RECT 0 28.035 0.070 28.385 ;
    RECT 0 28.455 0.070 28.805 ;
    RECT 0 28.875 0.070 29.225 ;
    RECT 0 29.295 0.070 29.645 ;
    RECT 0 29.715 0.070 31.885 ;
    RECT 0 31.955 0.070 32.305 ;
    RECT 0 32.375 0.070 32.725 ;
    RECT 0 32.795 0.070 33.145 ;
    RECT 0 33.215 0.070 33.565 ;
    RECT 0 33.635 0.070 33.985 ;
    RECT 0 34.055 0.070 34.405 ;
    RECT 0 34.475 0.070 34.825 ;
    RECT 0 34.895 0.070 35.245 ;
    RECT 0 35.315 0.070 35.665 ;
    RECT 0 35.735 0.070 36.085 ;
    RECT 0 36.155 0.070 36.505 ;
    RECT 0 36.575 0.070 36.925 ;
    RECT 0 36.995 0.070 37.345 ;
    RECT 0 37.415 0.070 37.765 ;
    RECT 0 37.835 0.070 38.185 ;
    RECT 0 38.255 0.070 38.605 ;
    RECT 0 38.675 0.070 39.025 ;
    RECT 0 39.095 0.070 39.445 ;
    RECT 0 39.515 0.070 39.865 ;
    RECT 0 39.935 0.070 40.285 ;
    RECT 0 40.355 0.070 40.705 ;
    RECT 0 40.775 0.070 41.125 ;
    RECT 0 41.195 0.070 41.545 ;
    RECT 0 41.615 0.070 41.965 ;
    RECT 0 42.035 0.070 42.385 ;
    RECT 0 42.455 0.070 42.805 ;
    RECT 0 42.875 0.070 43.225 ;
    RECT 0 43.295 0.070 43.645 ;
    RECT 0 43.715 0.070 44.065 ;
    RECT 0 44.135 0.070 44.485 ;
    RECT 0 44.555 0.070 44.905 ;
    RECT 0 44.975 0.070 47.145 ;
    RECT 0 47.215 0.070 47.565 ;
    RECT 0 47.635 0.070 47.985 ;
    RECT 0 48.055 0.070 48.405 ;
    RECT 0 48.475 0.070 48.825 ;
    RECT 0 48.895 0.070 49.245 ;
    RECT 0 49.315 0.070 51.485 ;
    RECT 0 51.555 0.070 51.905 ;
    RECT 0 51.975 0.070 52.325 ;
    RECT 0 52.395 0.070 56.000 ;
    LAYER metal4 ;
    RECT 0 0 19.190 1.400 ;
    RECT 0 54.600 19.190 56.000 ;
    RECT 0.000 1.400 1.260 54.600 ;
    RECT 1.540 1.400 2.380 54.600 ;
    RECT 2.660 1.400 3.500 54.600 ;
    RECT 3.780 1.400 4.620 54.600 ;
    RECT 4.900 1.400 5.740 54.600 ;
    RECT 6.020 1.400 6.860 54.600 ;
    RECT 7.140 1.400 7.980 54.600 ;
    RECT 8.260 1.400 9.100 54.600 ;
    RECT 9.380 1.400 10.220 54.600 ;
    RECT 10.500 1.400 11.340 54.600 ;
    RECT 11.620 1.400 12.460 54.600 ;
    RECT 12.740 1.400 13.580 54.600 ;
    RECT 13.860 1.400 14.700 54.600 ;
    RECT 14.980 1.400 15.820 54.600 ;
    RECT 16.100 1.400 16.940 54.600 ;
    RECT 17.220 1.400 19.190 54.600 ;
    LAYER via1 ;
    RECT 0 0 19.190 56.000 ;
    LAYER via2 ;
    RECT 0 0 19.190 56.000 ;
    LAYER via3 ;
    RECT 0 0 19.190 56.000 ;
    LAYER OVERLAP ;
    RECT 0 0 19.190 56.000 ;
  END
END fakeram45_64x32

END LIBRARY
